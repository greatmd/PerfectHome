# Created by MC2 : Version 2011.06.06 on 2013/09/17, 17:42:30

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2011.06.06
#        Technology     : 28 nm CMOS LOGIC High Performance Mobile 1P10M HKMG CU_ELK 0.9V
#        Memory Type    : TSMC 28nm High Performace Mobile Two Port Register File
#                       : with d240 bit cell Standard-Vt periphery
#        Library Name   : ts6n28hpma256x64m4f
#        Library Version: 110c
#        Generated Time : 2013/09/17, 17:42:29
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS6N28HPMA256X64M4F
	CLASS BLOCK ;
	FOREIGN TS6N28HPMA256X64M4F 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 47.765 BY 317.515 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 166.660 47.765 166.810 ;
			LAYER M3 ;
			RECT 47.525 166.660 47.765 166.810 ;
			LAYER M1 ;
			RECT 47.525 166.660 47.765 166.810 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 166.350 47.765 166.500 ;
			LAYER M1 ;
			RECT 47.525 166.350 47.765 166.500 ;
			LAYER M3 ;
			RECT 47.525 166.350 47.765 166.500 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 168.990 47.765 169.140 ;
			LAYER M2 ;
			RECT 47.525 168.990 47.765 169.140 ;
			LAYER M1 ;
			RECT 47.525 168.990 47.765 169.140 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 173.190 47.765 173.340 ;
			LAYER M2 ;
			RECT 47.525 173.190 47.765 173.340 ;
			LAYER M1 ;
			RECT 47.525 173.190 47.765 173.340 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[3]

	PIN AA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 170.240 47.765 170.390 ;
			LAYER M1 ;
			RECT 47.525 170.240 47.765 170.390 ;
			LAYER M2 ;
			RECT 47.525 170.240 47.765 170.390 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[4]

	PIN AA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 172.880 47.765 173.030 ;
			LAYER M2 ;
			RECT 47.525 172.880 47.765 173.030 ;
			LAYER M1 ;
			RECT 47.525 172.880 47.765 173.030 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[5]

	PIN AA[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 169.300 47.765 169.450 ;
			LAYER M3 ;
			RECT 47.525 169.300 47.765 169.450 ;
			LAYER M1 ;
			RECT 47.525 169.300 47.765 169.450 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[6]

	PIN AA[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 165.410 47.765 165.560 ;
			LAYER M2 ;
			RECT 47.525 165.410 47.765 165.560 ;
			LAYER M1 ;
			RECT 47.525 165.410 47.765 165.560 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AA[7]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 152.905 47.765 153.055 ;
			LAYER M1 ;
			RECT 47.525 152.905 47.765 153.055 ;
			LAYER M2 ;
			RECT 47.525 152.905 47.765 153.055 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 153.215 47.765 153.365 ;
			LAYER M2 ;
			RECT 47.525 153.215 47.765 153.365 ;
			LAYER M1 ;
			RECT 47.525 153.215 47.765 153.365 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 150.575 47.765 150.725 ;
			LAYER M1 ;
			RECT 47.525 150.575 47.765 150.725 ;
			LAYER M3 ;
			RECT 47.525 150.575 47.765 150.725 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.525 146.375 47.765 146.525 ;
			LAYER M3 ;
			RECT 47.525 146.375 47.765 146.525 ;
			LAYER M2 ;
			RECT 47.525 146.375 47.765 146.525 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[3]

	PIN AB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 149.325 47.765 149.475 ;
			LAYER M2 ;
			RECT 47.525 149.325 47.765 149.475 ;
			LAYER M1 ;
			RECT 47.525 149.325 47.765 149.475 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[4]

	PIN AB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 146.685 47.765 146.835 ;
			LAYER M3 ;
			RECT 47.525 146.685 47.765 146.835 ;
			LAYER M1 ;
			RECT 47.525 146.685 47.765 146.835 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[5]

	PIN AB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 150.265 47.765 150.415 ;
			LAYER M2 ;
			RECT 47.525 150.265 47.765 150.415 ;
			LAYER M1 ;
			RECT 47.525 150.265 47.765 150.415 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[6]

	PIN AB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.525 154.155 47.765 154.305 ;
			LAYER M3 ;
			RECT 47.525 154.155 47.765 154.305 ;
			LAYER M2 ;
			RECT 47.525 154.155 47.765 154.305 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0758 LAYER M1 ;
		ANTENNAMAXAREACAR 1.1371 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1575 LAYER M2 ;
		ANTENNAMAXAREACAR 5.6371 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 6.6657 LAYER M3 ;
	END AB[7]

	PIN CLKR
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 158.020 47.765 158.170 ;
			LAYER M2 ;
			RECT 47.525 158.020 47.765 158.170 ;
			LAYER M1 ;
			RECT 47.525 158.020 47.765 158.170 ;
		END
		ANTENNAGATEAREA 0.4767 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6122 LAYER M1 ;
		ANTENNAMAXAREACAR 6.7528 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0530 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4422 LAYER VIA1 ;
		ANTENNAGATEAREA 0.4767 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.3330 LAYER M2 ;
		ANTENNAMAXAREACAR 18.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.7755 LAYER VIA2 ;
		ANTENNAGATEAREA 0.4767 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.6379 LAYER M3 ;
		ANTENNAMAXAREACAR 19.7010 LAYER M3 ;
	END CLKR

	PIN CLKW
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 162.010 47.765 162.160 ;
			LAYER M2 ;
			RECT 47.525 162.010 47.765 162.160 ;
			LAYER M1 ;
			RECT 47.525 162.010 47.765 162.160 ;
		END
		ANTENNAGATEAREA 0.2185 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3678 LAYER M1 ;
		ANTENNAMAXAREACAR 9.4762 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0310 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.5159 LAYER VIA1 ;
		ANTENNAGATEAREA 0.2185 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.0483 LAYER M2 ;
		ANTENNAMAXAREACAR 18.0317 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0140 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8492 LAYER VIA2 ;
		ANTENNAGATEAREA 0.2185 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3566 LAYER M3 ;
		ANTENNAMAXAREACAR 19.6638 LAYER M3 ;
	END CLKW

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 3.715 47.765 3.955 ;
			LAYER M3 ;
			RECT 47.615 3.715 47.765 3.955 ;
			LAYER M2 ;
			RECT 47.615 3.715 47.765 3.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 47.715 47.765 47.955 ;
			LAYER M3 ;
			RECT 47.615 47.715 47.765 47.955 ;
			LAYER M1 ;
			RECT 47.615 47.715 47.765 47.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 52.115 47.765 52.355 ;
			LAYER M3 ;
			RECT 47.615 52.115 47.765 52.355 ;
			LAYER M1 ;
			RECT 47.615 52.115 47.765 52.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 56.515 47.765 56.755 ;
			LAYER M3 ;
			RECT 47.615 56.515 47.765 56.755 ;
			LAYER M1 ;
			RECT 47.615 56.515 47.765 56.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 60.915 47.765 61.155 ;
			LAYER M1 ;
			RECT 47.615 60.915 47.765 61.155 ;
			LAYER M3 ;
			RECT 47.615 60.915 47.765 61.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 65.315 47.765 65.555 ;
			LAYER M2 ;
			RECT 47.615 65.315 47.765 65.555 ;
			LAYER M3 ;
			RECT 47.615 65.315 47.765 65.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 69.715 47.765 69.955 ;
			LAYER M2 ;
			RECT 47.615 69.715 47.765 69.955 ;
			LAYER M3 ;
			RECT 47.615 69.715 47.765 69.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 74.115 47.765 74.355 ;
			LAYER M3 ;
			RECT 47.615 74.115 47.765 74.355 ;
			LAYER M2 ;
			RECT 47.615 74.115 47.765 74.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 78.515 47.765 78.755 ;
			LAYER M1 ;
			RECT 47.615 78.515 47.765 78.755 ;
			LAYER M3 ;
			RECT 47.615 78.515 47.765 78.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 82.915 47.765 83.155 ;
			LAYER M3 ;
			RECT 47.615 82.915 47.765 83.155 ;
			LAYER M2 ;
			RECT 47.615 82.915 47.765 83.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 87.315 47.765 87.555 ;
			LAYER M1 ;
			RECT 47.615 87.315 47.765 87.555 ;
			LAYER M3 ;
			RECT 47.615 87.315 47.765 87.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[19]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 8.115 47.765 8.355 ;
			LAYER M2 ;
			RECT 47.615 8.115 47.765 8.355 ;
			LAYER M1 ;
			RECT 47.615 8.115 47.765 8.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[1]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 91.715 47.765 91.955 ;
			LAYER M1 ;
			RECT 47.615 91.715 47.765 91.955 ;
			LAYER M3 ;
			RECT 47.615 91.715 47.765 91.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 96.115 47.765 96.355 ;
			LAYER M1 ;
			RECT 47.615 96.115 47.765 96.355 ;
			LAYER M3 ;
			RECT 47.615 96.115 47.765 96.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 100.515 47.765 100.755 ;
			LAYER M1 ;
			RECT 47.615 100.515 47.765 100.755 ;
			LAYER M3 ;
			RECT 47.615 100.515 47.765 100.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 104.915 47.765 105.155 ;
			LAYER M2 ;
			RECT 47.615 104.915 47.765 105.155 ;
			LAYER M1 ;
			RECT 47.615 104.915 47.765 105.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 109.315 47.765 109.555 ;
			LAYER M1 ;
			RECT 47.615 109.315 47.765 109.555 ;
			LAYER M3 ;
			RECT 47.615 109.315 47.765 109.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 113.715 47.765 113.955 ;
			LAYER M1 ;
			RECT 47.615 113.715 47.765 113.955 ;
			LAYER M2 ;
			RECT 47.615 113.715 47.765 113.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 118.115 47.765 118.355 ;
			LAYER M1 ;
			RECT 47.615 118.115 47.765 118.355 ;
			LAYER M3 ;
			RECT 47.615 118.115 47.765 118.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 122.515 47.765 122.755 ;
			LAYER M3 ;
			RECT 47.615 122.515 47.765 122.755 ;
			LAYER M2 ;
			RECT 47.615 122.515 47.765 122.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 126.915 47.765 127.155 ;
			LAYER M3 ;
			RECT 47.615 126.915 47.765 127.155 ;
			LAYER M2 ;
			RECT 47.615 126.915 47.765 127.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 131.315 47.765 131.555 ;
			LAYER M1 ;
			RECT 47.615 131.315 47.765 131.555 ;
			LAYER M2 ;
			RECT 47.615 131.315 47.765 131.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[29]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 12.515 47.765 12.755 ;
			LAYER M2 ;
			RECT 47.615 12.515 47.765 12.755 ;
			LAYER M1 ;
			RECT 47.615 12.515 47.765 12.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[2]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 135.715 47.765 135.955 ;
			LAYER M2 ;
			RECT 47.615 135.715 47.765 135.955 ;
			LAYER M1 ;
			RECT 47.615 135.715 47.765 135.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 140.115 47.765 140.355 ;
			LAYER M3 ;
			RECT 47.615 140.115 47.765 140.355 ;
			LAYER M1 ;
			RECT 47.615 140.115 47.765 140.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 178.730 47.765 178.970 ;
			LAYER M2 ;
			RECT 47.615 178.730 47.765 178.970 ;
			LAYER M1 ;
			RECT 47.615 178.730 47.765 178.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 183.130 47.765 183.370 ;
			LAYER M2 ;
			RECT 47.615 183.130 47.765 183.370 ;
			LAYER M3 ;
			RECT 47.615 183.130 47.765 183.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 187.530 47.765 187.770 ;
			LAYER M1 ;
			RECT 47.615 187.530 47.765 187.770 ;
			LAYER M2 ;
			RECT 47.615 187.530 47.765 187.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 191.930 47.765 192.170 ;
			LAYER M3 ;
			RECT 47.615 191.930 47.765 192.170 ;
			LAYER M2 ;
			RECT 47.615 191.930 47.765 192.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 196.330 47.765 196.570 ;
			LAYER M1 ;
			RECT 47.615 196.330 47.765 196.570 ;
			LAYER M2 ;
			RECT 47.615 196.330 47.765 196.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 200.730 47.765 200.970 ;
			LAYER M3 ;
			RECT 47.615 200.730 47.765 200.970 ;
			LAYER M2 ;
			RECT 47.615 200.730 47.765 200.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 205.130 47.765 205.370 ;
			LAYER M2 ;
			RECT 47.615 205.130 47.765 205.370 ;
			LAYER M1 ;
			RECT 47.615 205.130 47.765 205.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 209.530 47.765 209.770 ;
			LAYER M2 ;
			RECT 47.615 209.530 47.765 209.770 ;
			LAYER M1 ;
			RECT 47.615 209.530 47.765 209.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[39]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 16.915 47.765 17.155 ;
			LAYER M1 ;
			RECT 47.615 16.915 47.765 17.155 ;
			LAYER M3 ;
			RECT 47.615 16.915 47.765 17.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[3]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 213.930 47.765 214.170 ;
			LAYER M2 ;
			RECT 47.615 213.930 47.765 214.170 ;
			LAYER M3 ;
			RECT 47.615 213.930 47.765 214.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 218.330 47.765 218.570 ;
			LAYER M3 ;
			RECT 47.615 218.330 47.765 218.570 ;
			LAYER M2 ;
			RECT 47.615 218.330 47.765 218.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 222.730 47.765 222.970 ;
			LAYER M2 ;
			RECT 47.615 222.730 47.765 222.970 ;
			LAYER M1 ;
			RECT 47.615 222.730 47.765 222.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 227.130 47.765 227.370 ;
			LAYER M1 ;
			RECT 47.615 227.130 47.765 227.370 ;
			LAYER M3 ;
			RECT 47.615 227.130 47.765 227.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 231.530 47.765 231.770 ;
			LAYER M1 ;
			RECT 47.615 231.530 47.765 231.770 ;
			LAYER M3 ;
			RECT 47.615 231.530 47.765 231.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 235.930 47.765 236.170 ;
			LAYER M3 ;
			RECT 47.615 235.930 47.765 236.170 ;
			LAYER M2 ;
			RECT 47.615 235.930 47.765 236.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 240.330 47.765 240.570 ;
			LAYER M3 ;
			RECT 47.615 240.330 47.765 240.570 ;
			LAYER M2 ;
			RECT 47.615 240.330 47.765 240.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 244.730 47.765 244.970 ;
			LAYER M3 ;
			RECT 47.615 244.730 47.765 244.970 ;
			LAYER M1 ;
			RECT 47.615 244.730 47.765 244.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 249.130 47.765 249.370 ;
			LAYER M2 ;
			RECT 47.615 249.130 47.765 249.370 ;
			LAYER M1 ;
			RECT 47.615 249.130 47.765 249.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 253.530 47.765 253.770 ;
			LAYER M2 ;
			RECT 47.615 253.530 47.765 253.770 ;
			LAYER M3 ;
			RECT 47.615 253.530 47.765 253.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[49]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 21.315 47.765 21.555 ;
			LAYER M3 ;
			RECT 47.615 21.315 47.765 21.555 ;
			LAYER M2 ;
			RECT 47.615 21.315 47.765 21.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[4]

	PIN D[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 257.930 47.765 258.170 ;
			LAYER M2 ;
			RECT 47.615 257.930 47.765 258.170 ;
			LAYER M1 ;
			RECT 47.615 257.930 47.765 258.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[50]

	PIN D[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 262.330 47.765 262.570 ;
			LAYER M2 ;
			RECT 47.615 262.330 47.765 262.570 ;
			LAYER M3 ;
			RECT 47.615 262.330 47.765 262.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[51]

	PIN D[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 266.730 47.765 266.970 ;
			LAYER M2 ;
			RECT 47.615 266.730 47.765 266.970 ;
			LAYER M1 ;
			RECT 47.615 266.730 47.765 266.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[52]

	PIN D[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 271.130 47.765 271.370 ;
			LAYER M1 ;
			RECT 47.615 271.130 47.765 271.370 ;
			LAYER M2 ;
			RECT 47.615 271.130 47.765 271.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[53]

	PIN D[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 275.530 47.765 275.770 ;
			LAYER M1 ;
			RECT 47.615 275.530 47.765 275.770 ;
			LAYER M3 ;
			RECT 47.615 275.530 47.765 275.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[54]

	PIN D[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 279.930 47.765 280.170 ;
			LAYER M1 ;
			RECT 47.615 279.930 47.765 280.170 ;
			LAYER M3 ;
			RECT 47.615 279.930 47.765 280.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[55]

	PIN D[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 284.330 47.765 284.570 ;
			LAYER M1 ;
			RECT 47.615 284.330 47.765 284.570 ;
			LAYER M3 ;
			RECT 47.615 284.330 47.765 284.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[56]

	PIN D[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 288.730 47.765 288.970 ;
			LAYER M2 ;
			RECT 47.615 288.730 47.765 288.970 ;
			LAYER M1 ;
			RECT 47.615 288.730 47.765 288.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[57]

	PIN D[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 293.130 47.765 293.370 ;
			LAYER M2 ;
			RECT 47.615 293.130 47.765 293.370 ;
			LAYER M1 ;
			RECT 47.615 293.130 47.765 293.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[58]

	PIN D[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 297.530 47.765 297.770 ;
			LAYER M2 ;
			RECT 47.615 297.530 47.765 297.770 ;
			LAYER M1 ;
			RECT 47.615 297.530 47.765 297.770 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[59]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 25.715 47.765 25.955 ;
			LAYER M2 ;
			RECT 47.615 25.715 47.765 25.955 ;
			LAYER M3 ;
			RECT 47.615 25.715 47.765 25.955 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[5]

	PIN D[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 301.930 47.765 302.170 ;
			LAYER M3 ;
			RECT 47.615 301.930 47.765 302.170 ;
			LAYER M2 ;
			RECT 47.615 301.930 47.765 302.170 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[60]

	PIN D[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 306.330 47.765 306.570 ;
			LAYER M1 ;
			RECT 47.615 306.330 47.765 306.570 ;
			LAYER M3 ;
			RECT 47.615 306.330 47.765 306.570 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[61]

	PIN D[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 310.730 47.765 310.970 ;
			LAYER M3 ;
			RECT 47.615 310.730 47.765 310.970 ;
			LAYER M1 ;
			RECT 47.615 310.730 47.765 310.970 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[62]

	PIN D[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 315.130 47.765 315.370 ;
			LAYER M3 ;
			RECT 47.615 315.130 47.765 315.370 ;
			LAYER M1 ;
			RECT 47.615 315.130 47.765 315.370 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[63]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 30.115 47.765 30.355 ;
			LAYER M3 ;
			RECT 47.615 30.115 47.765 30.355 ;
			LAYER M2 ;
			RECT 47.615 30.115 47.765 30.355 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 34.515 47.765 34.755 ;
			LAYER M2 ;
			RECT 47.615 34.515 47.765 34.755 ;
			LAYER M1 ;
			RECT 47.615 34.515 47.765 34.755 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 38.915 47.765 39.155 ;
			LAYER M3 ;
			RECT 47.615 38.915 47.765 39.155 ;
			LAYER M2 ;
			RECT 47.615 38.915 47.765 39.155 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 43.315 47.765 43.555 ;
			LAYER M3 ;
			RECT 47.615 43.315 47.765 43.555 ;
			LAYER M2 ;
			RECT 47.615 43.315 47.765 43.555 ;
		END
		ANTENNAGATEAREA 0.0270 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.6796 LAYER M1 ;
		ANTENNAMAXAREACAR 2.2500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0220 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2407 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0270 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
		ANTENNAMAXAREACAR 8.3056 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4815 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0270 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 9.6389 LAYER M3 ;
	END D[9]

	PIN KP[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 155.335 47.765 155.485 ;
			LAYER M2 ;
			RECT 47.525 155.335 47.765 155.485 ;
			LAYER M1 ;
			RECT 47.525 155.335 47.765 155.485 ;
		END
		ANTENNAGATEAREA 0.1484 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3589 LAYER M1 ;
		ANTENNAMAXAREACAR 1.8302 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0330 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1348 LAYER VIA1 ;
		ANTENNAGATEAREA 0.1484 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 7.1721 LAYER M2 ;
		ANTENNAMAXAREACAR 63.6900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0310 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4852 LAYER VIA2 ;
		ANTENNAGATEAREA 0.1484 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5235 LAYER M3 ;
		ANTENNAMAXAREACAR 91.0755 LAYER M3 ;
	END KP[0]

	PIN KP[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 157.710 47.765 157.860 ;
			LAYER M3 ;
			RECT 47.525 157.710 47.765 157.860 ;
			LAYER M1 ;
			RECT 47.525 157.710 47.765 157.860 ;
		END
		ANTENNAGATEAREA 0.1484 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3589 LAYER M1 ;
		ANTENNAMAXAREACAR 1.8302 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0330 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1348 LAYER VIA1 ;
		ANTENNAGATEAREA 0.1484 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 7.1721 LAYER M2 ;
		ANTENNAMAXAREACAR 63.6900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0310 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4852 LAYER VIA2 ;
		ANTENNAGATEAREA 0.1484 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5235 LAYER M3 ;
		ANTENNAMAXAREACAR 91.0755 LAYER M3 ;
	END KP[1]

	PIN KP[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 157.090 47.765 157.240 ;
			LAYER M2 ;
			RECT 47.525 157.090 47.765 157.240 ;
			LAYER M1 ;
			RECT 47.525 157.090 47.765 157.240 ;
		END
		ANTENNAGATEAREA 0.1484 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3589 LAYER M1 ;
		ANTENNAMAXAREACAR 1.8302 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0330 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1348 LAYER VIA1 ;
		ANTENNAGATEAREA 0.1484 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 7.1721 LAYER M2 ;
		ANTENNAMAXAREACAR 63.6900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0310 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4852 LAYER VIA2 ;
		ANTENNAGATEAREA 0.1484 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5235 LAYER M3 ;
		ANTENNAMAXAREACAR 91.0755 LAYER M3 ;
	END KP[2]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 4.875 47.765 5.115 ;
			LAYER M2 ;
			RECT 47.615 4.875 47.765 5.115 ;
			LAYER M1 ;
			RECT 47.615 4.875 47.765 5.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 48.875 47.765 49.115 ;
			LAYER M3 ;
			RECT 47.615 48.875 47.765 49.115 ;
			LAYER M1 ;
			RECT 47.615 48.875 47.765 49.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 53.275 47.765 53.515 ;
			LAYER M1 ;
			RECT 47.615 53.275 47.765 53.515 ;
			LAYER M3 ;
			RECT 47.615 53.275 47.765 53.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 57.675 47.765 57.915 ;
			LAYER M3 ;
			RECT 47.615 57.675 47.765 57.915 ;
			LAYER M1 ;
			RECT 47.615 57.675 47.765 57.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 62.075 47.765 62.315 ;
			LAYER M3 ;
			RECT 47.615 62.075 47.765 62.315 ;
			LAYER M1 ;
			RECT 47.615 62.075 47.765 62.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 66.475 47.765 66.715 ;
			LAYER M1 ;
			RECT 47.615 66.475 47.765 66.715 ;
			LAYER M2 ;
			RECT 47.615 66.475 47.765 66.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 70.875 47.765 71.115 ;
			LAYER M2 ;
			RECT 47.615 70.875 47.765 71.115 ;
			LAYER M1 ;
			RECT 47.615 70.875 47.765 71.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 75.275 47.765 75.515 ;
			LAYER M1 ;
			RECT 47.615 75.275 47.765 75.515 ;
			LAYER M3 ;
			RECT 47.615 75.275 47.765 75.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 79.675 47.765 79.915 ;
			LAYER M3 ;
			RECT 47.615 79.675 47.765 79.915 ;
			LAYER M2 ;
			RECT 47.615 79.675 47.765 79.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 84.075 47.765 84.315 ;
			LAYER M3 ;
			RECT 47.615 84.075 47.765 84.315 ;
			LAYER M1 ;
			RECT 47.615 84.075 47.765 84.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 88.475 47.765 88.715 ;
			LAYER M2 ;
			RECT 47.615 88.475 47.765 88.715 ;
			LAYER M3 ;
			RECT 47.615 88.475 47.765 88.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[19]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 9.275 47.765 9.515 ;
			LAYER M3 ;
			RECT 47.615 9.275 47.765 9.515 ;
			LAYER M2 ;
			RECT 47.615 9.275 47.765 9.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[1]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 92.875 47.765 93.115 ;
			LAYER M2 ;
			RECT 47.615 92.875 47.765 93.115 ;
			LAYER M3 ;
			RECT 47.615 92.875 47.765 93.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 97.275 47.765 97.515 ;
			LAYER M3 ;
			RECT 47.615 97.275 47.765 97.515 ;
			LAYER M2 ;
			RECT 47.615 97.275 47.765 97.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 101.675 47.765 101.915 ;
			LAYER M2 ;
			RECT 47.615 101.675 47.765 101.915 ;
			LAYER M3 ;
			RECT 47.615 101.675 47.765 101.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 106.075 47.765 106.315 ;
			LAYER M3 ;
			RECT 47.615 106.075 47.765 106.315 ;
			LAYER M2 ;
			RECT 47.615 106.075 47.765 106.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 110.475 47.765 110.715 ;
			LAYER M1 ;
			RECT 47.615 110.475 47.765 110.715 ;
			LAYER M2 ;
			RECT 47.615 110.475 47.765 110.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 114.875 47.765 115.115 ;
			LAYER M2 ;
			RECT 47.615 114.875 47.765 115.115 ;
			LAYER M1 ;
			RECT 47.615 114.875 47.765 115.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 119.275 47.765 119.515 ;
			LAYER M1 ;
			RECT 47.615 119.275 47.765 119.515 ;
			LAYER M2 ;
			RECT 47.615 119.275 47.765 119.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 123.675 47.765 123.915 ;
			LAYER M2 ;
			RECT 47.615 123.675 47.765 123.915 ;
			LAYER M1 ;
			RECT 47.615 123.675 47.765 123.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 128.075 47.765 128.315 ;
			LAYER M3 ;
			RECT 47.615 128.075 47.765 128.315 ;
			LAYER M2 ;
			RECT 47.615 128.075 47.765 128.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 132.475 47.765 132.715 ;
			LAYER M3 ;
			RECT 47.615 132.475 47.765 132.715 ;
			LAYER M2 ;
			RECT 47.615 132.475 47.765 132.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[29]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 13.675 47.765 13.915 ;
			LAYER M3 ;
			RECT 47.615 13.675 47.765 13.915 ;
			LAYER M1 ;
			RECT 47.615 13.675 47.765 13.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[2]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 136.875 47.765 137.115 ;
			LAYER M3 ;
			RECT 47.615 136.875 47.765 137.115 ;
			LAYER M2 ;
			RECT 47.615 136.875 47.765 137.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 141.275 47.765 141.515 ;
			LAYER M1 ;
			RECT 47.615 141.275 47.765 141.515 ;
			LAYER M3 ;
			RECT 47.615 141.275 47.765 141.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 179.890 47.765 180.130 ;
			LAYER M3 ;
			RECT 47.615 179.890 47.765 180.130 ;
			LAYER M1 ;
			RECT 47.615 179.890 47.765 180.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 184.290 47.765 184.530 ;
			LAYER M3 ;
			RECT 47.615 184.290 47.765 184.530 ;
			LAYER M2 ;
			RECT 47.615 184.290 47.765 184.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 188.690 47.765 188.930 ;
			LAYER M2 ;
			RECT 47.615 188.690 47.765 188.930 ;
			LAYER M3 ;
			RECT 47.615 188.690 47.765 188.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 193.090 47.765 193.330 ;
			LAYER M3 ;
			RECT 47.615 193.090 47.765 193.330 ;
			LAYER M1 ;
			RECT 47.615 193.090 47.765 193.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 197.490 47.765 197.730 ;
			LAYER M1 ;
			RECT 47.615 197.490 47.765 197.730 ;
			LAYER M2 ;
			RECT 47.615 197.490 47.765 197.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 201.890 47.765 202.130 ;
			LAYER M2 ;
			RECT 47.615 201.890 47.765 202.130 ;
			LAYER M1 ;
			RECT 47.615 201.890 47.765 202.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 206.290 47.765 206.530 ;
			LAYER M1 ;
			RECT 47.615 206.290 47.765 206.530 ;
			LAYER M2 ;
			RECT 47.615 206.290 47.765 206.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 210.690 47.765 210.930 ;
			LAYER M2 ;
			RECT 47.615 210.690 47.765 210.930 ;
			LAYER M1 ;
			RECT 47.615 210.690 47.765 210.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[39]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 18.075 47.765 18.315 ;
			LAYER M2 ;
			RECT 47.615 18.075 47.765 18.315 ;
			LAYER M3 ;
			RECT 47.615 18.075 47.765 18.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[3]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 215.090 47.765 215.330 ;
			LAYER M1 ;
			RECT 47.615 215.090 47.765 215.330 ;
			LAYER M2 ;
			RECT 47.615 215.090 47.765 215.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 219.490 47.765 219.730 ;
			LAYER M3 ;
			RECT 47.615 219.490 47.765 219.730 ;
			LAYER M2 ;
			RECT 47.615 219.490 47.765 219.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 223.890 47.765 224.130 ;
			LAYER M2 ;
			RECT 47.615 223.890 47.765 224.130 ;
			LAYER M1 ;
			RECT 47.615 223.890 47.765 224.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 228.290 47.765 228.530 ;
			LAYER M2 ;
			RECT 47.615 228.290 47.765 228.530 ;
			LAYER M1 ;
			RECT 47.615 228.290 47.765 228.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 232.690 47.765 232.930 ;
			LAYER M2 ;
			RECT 47.615 232.690 47.765 232.930 ;
			LAYER M1 ;
			RECT 47.615 232.690 47.765 232.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 237.090 47.765 237.330 ;
			LAYER M1 ;
			RECT 47.615 237.090 47.765 237.330 ;
			LAYER M3 ;
			RECT 47.615 237.090 47.765 237.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 241.490 47.765 241.730 ;
			LAYER M2 ;
			RECT 47.615 241.490 47.765 241.730 ;
			LAYER M1 ;
			RECT 47.615 241.490 47.765 241.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 245.890 47.765 246.130 ;
			LAYER M1 ;
			RECT 47.615 245.890 47.765 246.130 ;
			LAYER M2 ;
			RECT 47.615 245.890 47.765 246.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 250.290 47.765 250.530 ;
			LAYER M3 ;
			RECT 47.615 250.290 47.765 250.530 ;
			LAYER M1 ;
			RECT 47.615 250.290 47.765 250.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 254.690 47.765 254.930 ;
			LAYER M2 ;
			RECT 47.615 254.690 47.765 254.930 ;
			LAYER M3 ;
			RECT 47.615 254.690 47.765 254.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[49]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 22.475 47.765 22.715 ;
			LAYER M3 ;
			RECT 47.615 22.475 47.765 22.715 ;
			LAYER M1 ;
			RECT 47.615 22.475 47.765 22.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[4]

	PIN Q[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 259.090 47.765 259.330 ;
			LAYER M2 ;
			RECT 47.615 259.090 47.765 259.330 ;
			LAYER M1 ;
			RECT 47.615 259.090 47.765 259.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[50]

	PIN Q[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 263.490 47.765 263.730 ;
			LAYER M2 ;
			RECT 47.615 263.490 47.765 263.730 ;
			LAYER M1 ;
			RECT 47.615 263.490 47.765 263.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[51]

	PIN Q[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 267.890 47.765 268.130 ;
			LAYER M2 ;
			RECT 47.615 267.890 47.765 268.130 ;
			LAYER M1 ;
			RECT 47.615 267.890 47.765 268.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[52]

	PIN Q[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 272.290 47.765 272.530 ;
			LAYER M1 ;
			RECT 47.615 272.290 47.765 272.530 ;
			LAYER M2 ;
			RECT 47.615 272.290 47.765 272.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[53]

	PIN Q[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 276.690 47.765 276.930 ;
			LAYER M3 ;
			RECT 47.615 276.690 47.765 276.930 ;
			LAYER M2 ;
			RECT 47.615 276.690 47.765 276.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[54]

	PIN Q[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 281.090 47.765 281.330 ;
			LAYER M2 ;
			RECT 47.615 281.090 47.765 281.330 ;
			LAYER M3 ;
			RECT 47.615 281.090 47.765 281.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[55]

	PIN Q[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 285.490 47.765 285.730 ;
			LAYER M3 ;
			RECT 47.615 285.490 47.765 285.730 ;
			LAYER M2 ;
			RECT 47.615 285.490 47.765 285.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[56]

	PIN Q[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 289.890 47.765 290.130 ;
			LAYER M3 ;
			RECT 47.615 289.890 47.765 290.130 ;
			LAYER M2 ;
			RECT 47.615 289.890 47.765 290.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[57]

	PIN Q[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 294.290 47.765 294.530 ;
			LAYER M1 ;
			RECT 47.615 294.290 47.765 294.530 ;
			LAYER M3 ;
			RECT 47.615 294.290 47.765 294.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[58]

	PIN Q[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 298.690 47.765 298.930 ;
			LAYER M2 ;
			RECT 47.615 298.690 47.765 298.930 ;
			LAYER M1 ;
			RECT 47.615 298.690 47.765 298.930 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[59]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 26.875 47.765 27.115 ;
			LAYER M1 ;
			RECT 47.615 26.875 47.765 27.115 ;
			LAYER M3 ;
			RECT 47.615 26.875 47.765 27.115 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[5]

	PIN Q[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 303.090 47.765 303.330 ;
			LAYER M1 ;
			RECT 47.615 303.090 47.765 303.330 ;
			LAYER M3 ;
			RECT 47.615 303.090 47.765 303.330 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[60]

	PIN Q[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 307.490 47.765 307.730 ;
			LAYER M2 ;
			RECT 47.615 307.490 47.765 307.730 ;
			LAYER M1 ;
			RECT 47.615 307.490 47.765 307.730 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[61]

	PIN Q[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 311.890 47.765 312.130 ;
			LAYER M1 ;
			RECT 47.615 311.890 47.765 312.130 ;
			LAYER M3 ;
			RECT 47.615 311.890 47.765 312.130 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[62]

	PIN Q[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.615 316.290 47.765 316.530 ;
			LAYER M1 ;
			RECT 47.615 316.290 47.765 316.530 ;
			LAYER M3 ;
			RECT 47.615 316.290 47.765 316.530 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[63]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 31.275 47.765 31.515 ;
			LAYER M2 ;
			RECT 47.615 31.275 47.765 31.515 ;
			LAYER M1 ;
			RECT 47.615 31.275 47.765 31.515 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 35.675 47.765 35.915 ;
			LAYER M2 ;
			RECT 47.615 35.675 47.765 35.915 ;
			LAYER M1 ;
			RECT 47.615 35.675 47.765 35.915 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.615 40.075 47.765 40.315 ;
			LAYER M2 ;
			RECT 47.615 40.075 47.765 40.315 ;
			LAYER M1 ;
			RECT 47.615 40.075 47.765 40.315 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.615 44.475 47.765 44.715 ;
			LAYER M2 ;
			RECT 47.615 44.475 47.765 44.715 ;
			LAYER M3 ;
			RECT 47.615 44.475 47.765 44.715 ;
		END
		ANTENNADIFFAREA 0.2120 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.3881 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0350 LAYER VIA1 ;
		ANTENNADIFFAREA 0.2120 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.5743 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNADIFFAREA 0.2120 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
	END Q[9]

	PIN RCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 151.505 47.765 151.655 ;
			LAYER M2 ;
			RECT 47.525 151.505 47.765 151.655 ;
			LAYER M1 ;
			RECT 47.525 151.505 47.765 151.655 ;
		END
		ANTENNAGATEAREA 0.0308 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1760 LAYER M1 ;
		ANTENNAMAXAREACAR 2.7922 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0280 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.3247 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0308 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.7790 LAYER M2 ;
		ANTENNAMAXAREACAR 28.0844 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0140 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.6169 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0308 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.1860 LAYER M3 ;
		ANTENNAMAXAREACAR 30.8117 LAYER M3 ;
	END RCT[0]

	PIN RCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.525 151.195 47.765 151.345 ;
			LAYER M3 ;
			RECT 47.525 151.195 47.765 151.345 ;
			LAYER M2 ;
			RECT 47.525 151.195 47.765 151.345 ;
		END
		ANTENNAGATEAREA 0.0308 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1760 LAYER M1 ;
		ANTENNAMAXAREACAR 2.7922 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0280 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.3247 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0308 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.7790 LAYER M2 ;
		ANTENNAMAXAREACAR 28.0844 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0140 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.6169 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0308 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.1860 LAYER M3 ;
		ANTENNAMAXAREACAR 30.8117 LAYER M3 ;
	END RCT[1]

	PIN REB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 155.955 47.765 156.105 ;
			LAYER M2 ;
			RECT 47.525 155.955 47.765 156.105 ;
			LAYER M1 ;
			RECT 47.525 155.955 47.765 156.105 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1953 LAYER M1 ;
		ANTENNAMAXAREACAR 4.5514 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0894 LAYER M2 ;
		ANTENNAMAXAREACAR 7.1057 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 8.1343 LAYER M3 ;
	END REB

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 1.805 47.765 2.095 ;
			LAYER M4 ;
			RECT 32.420 2.625 47.765 2.845 ;
			LAYER M4 ;
			RECT 0.000 4.005 47.765 4.295 ;
			LAYER M4 ;
			RECT 32.420 4.805 47.765 5.045 ;
			LAYER M4 ;
			RECT 0.000 6.205 47.765 6.495 ;
			LAYER M4 ;
			RECT 32.420 7.025 47.765 7.245 ;
			LAYER M4 ;
			RECT 0.000 8.405 47.765 8.695 ;
			LAYER M4 ;
			RECT 32.420 9.205 47.765 9.445 ;
			LAYER M4 ;
			RECT 0.000 10.605 47.765 10.895 ;
			LAYER M4 ;
			RECT 32.420 11.425 47.765 11.645 ;
			LAYER M4 ;
			RECT 0.000 12.805 47.765 13.095 ;
			LAYER M4 ;
			RECT 32.420 13.605 47.765 13.845 ;
			LAYER M4 ;
			RECT 0.000 15.005 47.765 15.295 ;
			LAYER M4 ;
			RECT 32.420 15.825 47.765 16.045 ;
			LAYER M4 ;
			RECT 0.000 17.205 47.765 17.495 ;
			LAYER M4 ;
			RECT 32.420 18.005 47.765 18.245 ;
			LAYER M4 ;
			RECT 0.000 19.405 47.765 19.695 ;
			LAYER M4 ;
			RECT 32.420 20.225 47.765 20.445 ;
			LAYER M4 ;
			RECT 0.000 21.605 47.765 21.895 ;
			LAYER M4 ;
			RECT 32.420 22.405 47.765 22.645 ;
			LAYER M4 ;
			RECT 0.000 23.805 47.765 24.095 ;
			LAYER M4 ;
			RECT 32.420 24.625 47.765 24.845 ;
			LAYER M4 ;
			RECT 0.000 26.005 47.765 26.295 ;
			LAYER M4 ;
			RECT 32.420 26.805 47.765 27.045 ;
			LAYER M4 ;
			RECT 0.000 28.205 47.765 28.495 ;
			LAYER M4 ;
			RECT 32.420 29.025 47.765 29.245 ;
			LAYER M4 ;
			RECT 0.000 30.405 47.765 30.695 ;
			LAYER M4 ;
			RECT 32.420 31.205 47.765 31.445 ;
			LAYER M4 ;
			RECT 0.000 32.605 47.765 32.895 ;
			LAYER M4 ;
			RECT 32.420 33.425 47.765 33.645 ;
			LAYER M4 ;
			RECT 0.000 34.805 47.765 35.095 ;
			LAYER M4 ;
			RECT 32.420 35.605 47.765 35.845 ;
			LAYER M4 ;
			RECT 0.000 37.005 47.765 37.295 ;
			LAYER M4 ;
			RECT 32.420 37.825 47.765 38.045 ;
			LAYER M4 ;
			RECT 0.000 39.205 47.765 39.495 ;
			LAYER M4 ;
			RECT 32.420 40.005 47.765 40.245 ;
			LAYER M4 ;
			RECT 0.000 41.405 47.765 41.695 ;
			LAYER M4 ;
			RECT 32.420 42.225 47.765 42.445 ;
			LAYER M4 ;
			RECT 0.000 43.605 47.765 43.895 ;
			LAYER M4 ;
			RECT 32.420 44.405 47.765 44.645 ;
			LAYER M4 ;
			RECT 0.000 45.805 47.765 46.095 ;
			LAYER M4 ;
			RECT 32.420 46.625 47.765 46.845 ;
			LAYER M4 ;
			RECT 0.000 48.005 47.765 48.295 ;
			LAYER M4 ;
			RECT 32.420 48.805 47.765 49.045 ;
			LAYER M4 ;
			RECT 0.000 50.205 47.765 50.495 ;
			LAYER M4 ;
			RECT 32.420 51.025 47.765 51.245 ;
			LAYER M4 ;
			RECT 0.000 52.405 47.765 52.695 ;
			LAYER M4 ;
			RECT 32.420 53.205 47.765 53.445 ;
			LAYER M4 ;
			RECT 0.000 54.605 47.765 54.895 ;
			LAYER M4 ;
			RECT 32.420 55.425 47.765 55.645 ;
			LAYER M4 ;
			RECT 0.000 56.805 47.765 57.095 ;
			LAYER M4 ;
			RECT 32.420 57.605 47.765 57.845 ;
			LAYER M4 ;
			RECT 0.000 59.005 47.765 59.295 ;
			LAYER M4 ;
			RECT 32.420 59.825 47.765 60.045 ;
			LAYER M4 ;
			RECT 0.000 61.205 47.765 61.495 ;
			LAYER M4 ;
			RECT 32.420 62.005 47.765 62.245 ;
			LAYER M4 ;
			RECT 0.000 63.405 47.765 63.695 ;
			LAYER M4 ;
			RECT 32.420 64.225 47.765 64.445 ;
			LAYER M4 ;
			RECT 0.000 65.605 47.765 65.895 ;
			LAYER M4 ;
			RECT 32.420 66.405 47.765 66.645 ;
			LAYER M4 ;
			RECT 0.000 67.805 47.765 68.095 ;
			LAYER M4 ;
			RECT 32.420 68.625 47.765 68.845 ;
			LAYER M4 ;
			RECT 0.000 70.005 47.765 70.295 ;
			LAYER M4 ;
			RECT 32.420 70.805 47.765 71.045 ;
			LAYER M4 ;
			RECT 0.000 72.205 47.765 72.495 ;
			LAYER M4 ;
			RECT 32.420 73.025 47.765 73.245 ;
			LAYER M4 ;
			RECT 0.000 74.405 47.765 74.695 ;
			LAYER M4 ;
			RECT 32.420 75.205 47.765 75.445 ;
			LAYER M4 ;
			RECT 0.000 76.605 47.765 76.895 ;
			LAYER M4 ;
			RECT 32.420 77.425 47.765 77.645 ;
			LAYER M4 ;
			RECT 0.000 78.805 47.765 79.095 ;
			LAYER M4 ;
			RECT 32.420 79.605 47.765 79.845 ;
			LAYER M4 ;
			RECT 0.000 81.005 47.765 81.295 ;
			LAYER M4 ;
			RECT 32.420 81.825 47.765 82.045 ;
			LAYER M4 ;
			RECT 0.000 83.205 47.765 83.495 ;
			LAYER M4 ;
			RECT 32.420 84.005 47.765 84.245 ;
			LAYER M4 ;
			RECT 0.000 85.405 47.765 85.695 ;
			LAYER M4 ;
			RECT 32.420 86.225 47.765 86.445 ;
			LAYER M4 ;
			RECT 0.000 87.605 47.765 87.895 ;
			LAYER M4 ;
			RECT 32.420 88.405 47.765 88.645 ;
			LAYER M4 ;
			RECT 0.000 89.805 47.765 90.095 ;
			LAYER M4 ;
			RECT 32.420 90.625 47.765 90.845 ;
			LAYER M4 ;
			RECT 0.000 92.005 47.765 92.295 ;
			LAYER M4 ;
			RECT 32.420 92.805 47.765 93.045 ;
			LAYER M4 ;
			RECT 0.000 94.205 47.765 94.495 ;
			LAYER M4 ;
			RECT 32.420 95.025 47.765 95.245 ;
			LAYER M4 ;
			RECT 0.000 96.405 47.765 96.695 ;
			LAYER M4 ;
			RECT 32.420 97.205 47.765 97.445 ;
			LAYER M4 ;
			RECT 0.000 98.605 47.765 98.895 ;
			LAYER M4 ;
			RECT 32.420 99.425 47.765 99.645 ;
			LAYER M4 ;
			RECT 0.000 100.805 47.765 101.095 ;
			LAYER M4 ;
			RECT 32.420 101.605 47.765 101.845 ;
			LAYER M4 ;
			RECT 0.000 103.005 47.765 103.295 ;
			LAYER M4 ;
			RECT 32.420 103.825 47.765 104.045 ;
			LAYER M4 ;
			RECT 0.000 105.205 47.765 105.495 ;
			LAYER M4 ;
			RECT 32.420 106.005 47.765 106.245 ;
			LAYER M4 ;
			RECT 0.000 107.405 47.765 107.695 ;
			LAYER M4 ;
			RECT 32.420 108.225 47.765 108.445 ;
			LAYER M4 ;
			RECT 0.000 109.605 47.765 109.895 ;
			LAYER M4 ;
			RECT 32.420 110.405 47.765 110.645 ;
			LAYER M4 ;
			RECT 0.000 111.805 47.765 112.095 ;
			LAYER M4 ;
			RECT 32.420 112.625 47.765 112.845 ;
			LAYER M4 ;
			RECT 0.000 114.005 47.765 114.295 ;
			LAYER M4 ;
			RECT 32.420 114.805 47.765 115.045 ;
			LAYER M4 ;
			RECT 0.000 116.205 47.765 116.495 ;
			LAYER M4 ;
			RECT 32.420 117.025 47.765 117.245 ;
			LAYER M4 ;
			RECT 0.000 118.405 47.765 118.695 ;
			LAYER M4 ;
			RECT 32.420 119.205 47.765 119.445 ;
			LAYER M4 ;
			RECT 0.000 120.605 47.765 120.895 ;
			LAYER M4 ;
			RECT 32.420 121.425 47.765 121.645 ;
			LAYER M4 ;
			RECT 0.000 122.805 47.765 123.095 ;
			LAYER M4 ;
			RECT 32.420 123.605 47.765 123.845 ;
			LAYER M4 ;
			RECT 0.000 125.005 47.765 125.295 ;
			LAYER M4 ;
			RECT 32.420 125.825 47.765 126.045 ;
			LAYER M4 ;
			RECT 0.000 127.205 47.765 127.495 ;
			LAYER M4 ;
			RECT 32.420 128.005 47.765 128.245 ;
			LAYER M4 ;
			RECT 0.000 129.405 47.765 129.695 ;
			LAYER M4 ;
			RECT 32.420 130.225 47.765 130.445 ;
			LAYER M4 ;
			RECT 0.000 131.605 47.765 131.895 ;
			LAYER M4 ;
			RECT 32.420 132.405 47.765 132.645 ;
			LAYER M4 ;
			RECT 0.000 133.805 47.765 134.095 ;
			LAYER M4 ;
			RECT 32.420 134.625 47.765 134.845 ;
			LAYER M4 ;
			RECT 0.000 136.005 47.765 136.295 ;
			LAYER M4 ;
			RECT 32.420 136.805 47.765 137.045 ;
			LAYER M4 ;
			RECT 0.000 138.205 47.765 138.495 ;
			LAYER M4 ;
			RECT 32.420 139.025 47.765 139.245 ;
			LAYER M4 ;
			RECT 0.000 140.405 47.765 140.695 ;
			LAYER M4 ;
			RECT 32.420 141.205 47.765 141.445 ;
			LAYER M4 ;
			RECT 32.420 141.855 47.765 142.095 ;
			LAYER M4 ;
			RECT 0.000 142.605 47.765 142.895 ;
			LAYER M4 ;
			RECT 0.000 147.270 47.765 147.770 ;
			LAYER M4 ;
			RECT 0.000 150.670 47.765 151.270 ;
			LAYER M4 ;
			RECT 0.000 152.580 47.765 153.180 ;
			LAYER M4 ;
			RECT 0.000 155.520 47.765 155.970 ;
			LAYER M4 ;
			RECT 0.000 158.280 47.765 158.730 ;
			LAYER M4 ;
			RECT 0.000 161.070 47.765 161.670 ;
			LAYER M4 ;
			RECT 0.000 162.980 47.765 163.580 ;
			LAYER M4 ;
			RECT 0.000 166.480 47.765 166.980 ;
			LAYER M4 ;
			RECT 0.000 174.620 47.765 174.910 ;
			LAYER M4 ;
			RECT 32.420 175.420 47.765 175.660 ;
			LAYER M4 ;
			RECT 0.000 176.820 47.765 177.110 ;
			LAYER M4 ;
			RECT 32.420 177.640 47.765 177.860 ;
			LAYER M4 ;
			RECT 0.000 179.020 47.765 179.310 ;
			LAYER M4 ;
			RECT 32.420 179.820 47.765 180.060 ;
			LAYER M4 ;
			RECT 0.000 181.220 47.765 181.510 ;
			LAYER M4 ;
			RECT 32.420 182.040 47.765 182.260 ;
			LAYER M4 ;
			RECT 0.000 183.420 47.765 183.710 ;
			LAYER M4 ;
			RECT 32.420 184.220 47.765 184.460 ;
			LAYER M4 ;
			RECT 0.000 185.620 47.765 185.910 ;
			LAYER M4 ;
			RECT 32.420 186.440 47.765 186.660 ;
			LAYER M4 ;
			RECT 0.000 187.820 47.765 188.110 ;
			LAYER M4 ;
			RECT 32.420 188.620 47.765 188.860 ;
			LAYER M4 ;
			RECT 0.000 190.020 47.765 190.310 ;
			LAYER M4 ;
			RECT 32.420 190.840 47.765 191.060 ;
			LAYER M4 ;
			RECT 0.000 192.220 47.765 192.510 ;
			LAYER M4 ;
			RECT 32.420 193.020 47.765 193.260 ;
			LAYER M4 ;
			RECT 0.000 194.420 47.765 194.710 ;
			LAYER M4 ;
			RECT 32.420 195.240 47.765 195.460 ;
			LAYER M4 ;
			RECT 0.000 196.620 47.765 196.910 ;
			LAYER M4 ;
			RECT 32.420 197.420 47.765 197.660 ;
			LAYER M4 ;
			RECT 0.000 198.820 47.765 199.110 ;
			LAYER M4 ;
			RECT 32.420 199.640 47.765 199.860 ;
			LAYER M4 ;
			RECT 0.000 201.020 47.765 201.310 ;
			LAYER M4 ;
			RECT 32.420 201.820 47.765 202.060 ;
			LAYER M4 ;
			RECT 0.000 203.220 47.765 203.510 ;
			LAYER M4 ;
			RECT 32.420 204.040 47.765 204.260 ;
			LAYER M4 ;
			RECT 0.000 205.420 47.765 205.710 ;
			LAYER M4 ;
			RECT 32.420 206.220 47.765 206.460 ;
			LAYER M4 ;
			RECT 0.000 207.620 47.765 207.910 ;
			LAYER M4 ;
			RECT 32.420 208.440 47.765 208.660 ;
			LAYER M4 ;
			RECT 0.000 209.820 47.765 210.110 ;
			LAYER M4 ;
			RECT 32.420 210.620 47.765 210.860 ;
			LAYER M4 ;
			RECT 0.000 212.020 47.765 212.310 ;
			LAYER M4 ;
			RECT 32.420 212.840 47.765 213.060 ;
			LAYER M4 ;
			RECT 0.000 214.220 47.765 214.510 ;
			LAYER M4 ;
			RECT 32.420 215.020 47.765 215.260 ;
			LAYER M4 ;
			RECT 0.000 216.420 47.765 216.710 ;
			LAYER M4 ;
			RECT 32.420 217.240 47.765 217.460 ;
			LAYER M4 ;
			RECT 0.000 218.620 47.765 218.910 ;
			LAYER M4 ;
			RECT 32.420 219.420 47.765 219.660 ;
			LAYER M4 ;
			RECT 0.000 220.820 47.765 221.110 ;
			LAYER M4 ;
			RECT 32.420 221.640 47.765 221.860 ;
			LAYER M4 ;
			RECT 0.000 223.020 47.765 223.310 ;
			LAYER M4 ;
			RECT 32.420 223.820 47.765 224.060 ;
			LAYER M4 ;
			RECT 0.000 225.220 47.765 225.510 ;
			LAYER M4 ;
			RECT 32.420 226.040 47.765 226.260 ;
			LAYER M4 ;
			RECT 0.000 227.420 47.765 227.710 ;
			LAYER M4 ;
			RECT 32.420 228.220 47.765 228.460 ;
			LAYER M4 ;
			RECT 0.000 229.620 47.765 229.910 ;
			LAYER M4 ;
			RECT 32.420 230.440 47.765 230.660 ;
			LAYER M4 ;
			RECT 0.000 231.820 47.765 232.110 ;
			LAYER M4 ;
			RECT 32.420 232.620 47.765 232.860 ;
			LAYER M4 ;
			RECT 0.000 234.020 47.765 234.310 ;
			LAYER M4 ;
			RECT 32.420 234.840 47.765 235.060 ;
			LAYER M4 ;
			RECT 0.000 236.220 47.765 236.510 ;
			LAYER M4 ;
			RECT 32.420 237.020 47.765 237.260 ;
			LAYER M4 ;
			RECT 0.000 238.420 47.765 238.710 ;
			LAYER M4 ;
			RECT 32.420 239.240 47.765 239.460 ;
			LAYER M4 ;
			RECT 0.000 240.620 47.765 240.910 ;
			LAYER M4 ;
			RECT 32.420 241.420 47.765 241.660 ;
			LAYER M4 ;
			RECT 0.000 242.820 47.765 243.110 ;
			LAYER M4 ;
			RECT 32.420 243.640 47.765 243.860 ;
			LAYER M4 ;
			RECT 0.000 245.020 47.765 245.310 ;
			LAYER M4 ;
			RECT 32.420 245.820 47.765 246.060 ;
			LAYER M4 ;
			RECT 0.000 247.220 47.765 247.510 ;
			LAYER M4 ;
			RECT 32.420 248.040 47.765 248.260 ;
			LAYER M4 ;
			RECT 0.000 249.420 47.765 249.710 ;
			LAYER M4 ;
			RECT 32.420 250.220 47.765 250.460 ;
			LAYER M4 ;
			RECT 0.000 251.620 47.765 251.910 ;
			LAYER M4 ;
			RECT 32.420 252.440 47.765 252.660 ;
			LAYER M4 ;
			RECT 0.000 253.820 47.765 254.110 ;
			LAYER M4 ;
			RECT 32.420 254.620 47.765 254.860 ;
			LAYER M4 ;
			RECT 0.000 256.020 47.765 256.310 ;
			LAYER M4 ;
			RECT 32.420 256.840 47.765 257.060 ;
			LAYER M4 ;
			RECT 0.000 258.220 47.765 258.510 ;
			LAYER M4 ;
			RECT 32.420 259.020 47.765 259.260 ;
			LAYER M4 ;
			RECT 0.000 260.420 47.765 260.710 ;
			LAYER M4 ;
			RECT 32.420 261.240 47.765 261.460 ;
			LAYER M4 ;
			RECT 0.000 262.620 47.765 262.910 ;
			LAYER M4 ;
			RECT 32.420 263.420 47.765 263.660 ;
			LAYER M4 ;
			RECT 0.000 264.820 47.765 265.110 ;
			LAYER M4 ;
			RECT 32.420 265.640 47.765 265.860 ;
			LAYER M4 ;
			RECT 0.000 267.020 47.765 267.310 ;
			LAYER M4 ;
			RECT 32.420 267.820 47.765 268.060 ;
			LAYER M4 ;
			RECT 0.000 269.220 47.765 269.510 ;
			LAYER M4 ;
			RECT 32.420 270.040 47.765 270.260 ;
			LAYER M4 ;
			RECT 0.000 271.420 47.765 271.710 ;
			LAYER M4 ;
			RECT 32.420 272.220 47.765 272.460 ;
			LAYER M4 ;
			RECT 0.000 273.620 47.765 273.910 ;
			LAYER M4 ;
			RECT 32.420 274.440 47.765 274.660 ;
			LAYER M4 ;
			RECT 0.000 275.820 47.765 276.110 ;
			LAYER M4 ;
			RECT 32.420 276.620 47.765 276.860 ;
			LAYER M4 ;
			RECT 0.000 278.020 47.765 278.310 ;
			LAYER M4 ;
			RECT 32.420 278.840 47.765 279.060 ;
			LAYER M4 ;
			RECT 0.000 280.220 47.765 280.510 ;
			LAYER M4 ;
			RECT 32.420 281.020 47.765 281.260 ;
			LAYER M4 ;
			RECT 0.000 282.420 47.765 282.710 ;
			LAYER M4 ;
			RECT 32.420 283.240 47.765 283.460 ;
			LAYER M4 ;
			RECT 0.000 284.620 47.765 284.910 ;
			LAYER M4 ;
			RECT 32.420 285.420 47.765 285.660 ;
			LAYER M4 ;
			RECT 0.000 286.820 47.765 287.110 ;
			LAYER M4 ;
			RECT 32.420 287.640 47.765 287.860 ;
			LAYER M4 ;
			RECT 0.000 289.020 47.765 289.310 ;
			LAYER M4 ;
			RECT 32.420 289.820 47.765 290.060 ;
			LAYER M4 ;
			RECT 0.000 291.220 47.765 291.510 ;
			LAYER M4 ;
			RECT 32.420 292.040 47.765 292.260 ;
			LAYER M4 ;
			RECT 0.000 293.420 47.765 293.710 ;
			LAYER M4 ;
			RECT 32.420 294.220 47.765 294.460 ;
			LAYER M4 ;
			RECT 0.000 295.620 47.765 295.910 ;
			LAYER M4 ;
			RECT 32.420 296.440 47.765 296.660 ;
			LAYER M4 ;
			RECT 0.000 297.820 47.765 298.110 ;
			LAYER M4 ;
			RECT 32.420 298.620 47.765 298.860 ;
			LAYER M4 ;
			RECT 0.000 300.020 47.765 300.310 ;
			LAYER M4 ;
			RECT 32.420 300.840 47.765 301.060 ;
			LAYER M4 ;
			RECT 0.000 302.220 47.765 302.510 ;
			LAYER M4 ;
			RECT 32.420 303.020 47.765 303.260 ;
			LAYER M4 ;
			RECT 0.000 304.420 47.765 304.710 ;
			LAYER M4 ;
			RECT 32.420 305.240 47.765 305.460 ;
			LAYER M4 ;
			RECT 0.000 306.620 47.765 306.910 ;
			LAYER M4 ;
			RECT 32.420 307.420 47.765 307.660 ;
			LAYER M4 ;
			RECT 0.000 308.820 47.765 309.110 ;
			LAYER M4 ;
			RECT 32.420 309.640 47.765 309.860 ;
			LAYER M4 ;
			RECT 0.000 311.020 47.765 311.310 ;
			LAYER M4 ;
			RECT 32.420 311.820 47.765 312.060 ;
			LAYER M4 ;
			RECT 0.000 313.220 47.765 313.510 ;
			LAYER M4 ;
			RECT 32.420 314.040 47.765 314.260 ;
			LAYER M4 ;
			RECT 0.000 315.420 47.765 315.710 ;
			LAYER M4 ;
			RECT 32.420 316.220 47.765 316.460 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 0.745 47.765 0.955 ;
			LAYER M4 ;
			RECT 32.420 1.055 47.765 1.295 ;
			LAYER M4 ;
			RECT 0.000 2.945 47.765 3.155 ;
			LAYER M4 ;
			RECT 32.420 3.255 47.765 3.475 ;
			LAYER M4 ;
			RECT 0.000 5.145 47.765 5.355 ;
			LAYER M4 ;
			RECT 32.420 5.455 47.765 5.695 ;
			LAYER M4 ;
			RECT 0.000 7.345 47.765 7.555 ;
			LAYER M4 ;
			RECT 32.420 7.655 47.765 7.875 ;
			LAYER M4 ;
			RECT 0.000 9.545 47.765 9.755 ;
			LAYER M4 ;
			RECT 32.420 9.855 47.765 10.095 ;
			LAYER M4 ;
			RECT 0.000 11.745 47.765 11.955 ;
			LAYER M4 ;
			RECT 32.420 12.055 47.765 12.275 ;
			LAYER M4 ;
			RECT 0.000 13.945 47.765 14.155 ;
			LAYER M4 ;
			RECT 32.420 14.255 47.765 14.495 ;
			LAYER M4 ;
			RECT 0.000 16.145 47.765 16.355 ;
			LAYER M4 ;
			RECT 32.420 16.455 47.765 16.675 ;
			LAYER M4 ;
			RECT 0.000 18.345 47.765 18.555 ;
			LAYER M4 ;
			RECT 32.420 18.655 47.765 18.895 ;
			LAYER M4 ;
			RECT 0.000 20.545 47.765 20.755 ;
			LAYER M4 ;
			RECT 32.420 20.855 47.765 21.075 ;
			LAYER M4 ;
			RECT 0.000 22.745 47.765 22.955 ;
			LAYER M4 ;
			RECT 32.420 23.055 47.765 23.295 ;
			LAYER M4 ;
			RECT 0.000 24.945 47.765 25.155 ;
			LAYER M4 ;
			RECT 32.420 25.255 47.765 25.475 ;
			LAYER M4 ;
			RECT 0.000 27.145 47.765 27.355 ;
			LAYER M4 ;
			RECT 32.420 27.455 47.765 27.695 ;
			LAYER M4 ;
			RECT 0.000 29.345 47.765 29.555 ;
			LAYER M4 ;
			RECT 32.420 29.655 47.765 29.875 ;
			LAYER M4 ;
			RECT 0.000 31.545 47.765 31.755 ;
			LAYER M4 ;
			RECT 32.420 31.855 47.765 32.095 ;
			LAYER M4 ;
			RECT 0.000 33.745 47.765 33.955 ;
			LAYER M4 ;
			RECT 32.420 34.055 47.765 34.275 ;
			LAYER M4 ;
			RECT 0.000 35.945 47.765 36.155 ;
			LAYER M4 ;
			RECT 32.420 36.255 47.765 36.495 ;
			LAYER M4 ;
			RECT 0.000 38.145 47.765 38.355 ;
			LAYER M4 ;
			RECT 32.420 38.455 47.765 38.675 ;
			LAYER M4 ;
			RECT 0.000 40.345 47.765 40.555 ;
			LAYER M4 ;
			RECT 32.420 40.655 47.765 40.895 ;
			LAYER M4 ;
			RECT 0.000 42.545 47.765 42.755 ;
			LAYER M4 ;
			RECT 32.420 42.855 47.765 43.075 ;
			LAYER M4 ;
			RECT 0.000 44.745 47.765 44.955 ;
			LAYER M4 ;
			RECT 32.420 45.055 47.765 45.295 ;
			LAYER M4 ;
			RECT 0.000 46.945 47.765 47.155 ;
			LAYER M4 ;
			RECT 32.420 47.255 47.765 47.475 ;
			LAYER M4 ;
			RECT 0.000 49.145 47.765 49.355 ;
			LAYER M4 ;
			RECT 32.420 49.455 47.765 49.695 ;
			LAYER M4 ;
			RECT 0.000 51.345 47.765 51.555 ;
			LAYER M4 ;
			RECT 32.420 51.655 47.765 51.875 ;
			LAYER M4 ;
			RECT 0.000 53.545 47.765 53.755 ;
			LAYER M4 ;
			RECT 32.420 53.855 47.765 54.095 ;
			LAYER M4 ;
			RECT 0.000 55.745 47.765 55.955 ;
			LAYER M4 ;
			RECT 32.420 56.055 47.765 56.275 ;
			LAYER M4 ;
			RECT 0.000 57.945 47.765 58.155 ;
			LAYER M4 ;
			RECT 32.420 58.255 47.765 58.495 ;
			LAYER M4 ;
			RECT 0.000 60.145 47.765 60.355 ;
			LAYER M4 ;
			RECT 32.420 60.455 47.765 60.675 ;
			LAYER M4 ;
			RECT 0.000 62.345 47.765 62.555 ;
			LAYER M4 ;
			RECT 32.420 62.655 47.765 62.895 ;
			LAYER M4 ;
			RECT 0.000 64.545 47.765 64.755 ;
			LAYER M4 ;
			RECT 32.420 64.855 47.765 65.075 ;
			LAYER M4 ;
			RECT 0.000 66.745 47.765 66.955 ;
			LAYER M4 ;
			RECT 32.420 67.055 47.765 67.295 ;
			LAYER M4 ;
			RECT 0.000 68.945 47.765 69.155 ;
			LAYER M4 ;
			RECT 32.420 69.255 47.765 69.475 ;
			LAYER M4 ;
			RECT 0.000 71.145 47.765 71.355 ;
			LAYER M4 ;
			RECT 32.420 71.455 47.765 71.695 ;
			LAYER M4 ;
			RECT 0.000 73.345 47.765 73.555 ;
			LAYER M4 ;
			RECT 32.420 73.655 47.765 73.875 ;
			LAYER M4 ;
			RECT 0.000 75.545 47.765 75.755 ;
			LAYER M4 ;
			RECT 32.420 75.855 47.765 76.095 ;
			LAYER M4 ;
			RECT 0.000 77.745 47.765 77.955 ;
			LAYER M4 ;
			RECT 32.420 78.055 47.765 78.275 ;
			LAYER M4 ;
			RECT 0.000 79.945 47.765 80.155 ;
			LAYER M4 ;
			RECT 32.420 80.255 47.765 80.495 ;
			LAYER M4 ;
			RECT 0.000 82.145 47.765 82.355 ;
			LAYER M4 ;
			RECT 32.420 82.455 47.765 82.675 ;
			LAYER M4 ;
			RECT 0.000 84.345 47.765 84.555 ;
			LAYER M4 ;
			RECT 32.420 84.655 47.765 84.895 ;
			LAYER M4 ;
			RECT 0.000 86.545 47.765 86.755 ;
			LAYER M4 ;
			RECT 32.420 86.855 47.765 87.075 ;
			LAYER M4 ;
			RECT 0.000 88.745 47.765 88.955 ;
			LAYER M4 ;
			RECT 32.420 89.055 47.765 89.295 ;
			LAYER M4 ;
			RECT 0.000 90.945 47.765 91.155 ;
			LAYER M4 ;
			RECT 32.420 91.255 47.765 91.475 ;
			LAYER M4 ;
			RECT 0.000 93.145 47.765 93.355 ;
			LAYER M4 ;
			RECT 32.420 93.455 47.765 93.695 ;
			LAYER M4 ;
			RECT 0.000 95.345 47.765 95.555 ;
			LAYER M4 ;
			RECT 32.420 95.655 47.765 95.875 ;
			LAYER M4 ;
			RECT 0.000 97.545 47.765 97.755 ;
			LAYER M4 ;
			RECT 32.420 97.855 47.765 98.095 ;
			LAYER M4 ;
			RECT 0.000 99.745 47.765 99.955 ;
			LAYER M4 ;
			RECT 32.420 100.055 47.765 100.275 ;
			LAYER M4 ;
			RECT 0.000 101.945 47.765 102.155 ;
			LAYER M4 ;
			RECT 32.420 102.255 47.765 102.495 ;
			LAYER M4 ;
			RECT 0.000 104.145 47.765 104.355 ;
			LAYER M4 ;
			RECT 32.420 104.455 47.765 104.675 ;
			LAYER M4 ;
			RECT 0.000 106.345 47.765 106.555 ;
			LAYER M4 ;
			RECT 32.420 106.655 47.765 106.895 ;
			LAYER M4 ;
			RECT 0.000 108.545 47.765 108.755 ;
			LAYER M4 ;
			RECT 32.420 108.855 47.765 109.075 ;
			LAYER M4 ;
			RECT 0.000 110.745 47.765 110.955 ;
			LAYER M4 ;
			RECT 32.420 111.055 47.765 111.295 ;
			LAYER M4 ;
			RECT 0.000 112.945 47.765 113.155 ;
			LAYER M4 ;
			RECT 32.420 113.255 47.765 113.475 ;
			LAYER M4 ;
			RECT 0.000 115.145 47.765 115.355 ;
			LAYER M4 ;
			RECT 32.420 115.455 47.765 115.695 ;
			LAYER M4 ;
			RECT 0.000 117.345 47.765 117.555 ;
			LAYER M4 ;
			RECT 32.420 117.655 47.765 117.875 ;
			LAYER M4 ;
			RECT 0.000 119.545 47.765 119.755 ;
			LAYER M4 ;
			RECT 32.420 119.855 47.765 120.095 ;
			LAYER M4 ;
			RECT 0.000 121.745 47.765 121.955 ;
			LAYER M4 ;
			RECT 32.420 122.055 47.765 122.275 ;
			LAYER M4 ;
			RECT 0.000 123.945 47.765 124.155 ;
			LAYER M4 ;
			RECT 32.420 124.255 47.765 124.495 ;
			LAYER M4 ;
			RECT 0.000 126.145 47.765 126.355 ;
			LAYER M4 ;
			RECT 32.420 126.455 47.765 126.675 ;
			LAYER M4 ;
			RECT 0.000 128.345 47.765 128.555 ;
			LAYER M4 ;
			RECT 32.420 128.655 47.765 128.895 ;
			LAYER M4 ;
			RECT 0.000 130.545 47.765 130.755 ;
			LAYER M4 ;
			RECT 32.420 130.855 47.765 131.075 ;
			LAYER M4 ;
			RECT 0.000 132.745 47.765 132.955 ;
			LAYER M4 ;
			RECT 32.420 133.055 47.765 133.295 ;
			LAYER M4 ;
			RECT 0.000 134.945 47.765 135.155 ;
			LAYER M4 ;
			RECT 32.420 135.255 47.765 135.475 ;
			LAYER M4 ;
			RECT 0.000 137.145 47.765 137.355 ;
			LAYER M4 ;
			RECT 32.420 137.455 47.765 137.695 ;
			LAYER M4 ;
			RECT 0.000 139.345 47.765 139.555 ;
			LAYER M4 ;
			RECT 32.420 139.655 47.765 139.875 ;
			LAYER M4 ;
			RECT 0.000 141.545 47.765 141.755 ;
			LAYER M4 ;
			RECT 32.420 143.405 47.765 143.645 ;
			LAYER M4 ;
			RECT 0.000 143.745 47.765 143.955 ;
			LAYER M4 ;
			RECT 0.000 144.300 47.765 144.700 ;
			LAYER M4 ;
			RECT 0.000 144.830 47.765 145.330 ;
			LAYER M4 ;
			RECT 0.000 146.640 47.765 147.140 ;
			LAYER M4 ;
			RECT 0.000 148.530 47.765 149.030 ;
			LAYER M4 ;
			RECT 0.000 153.310 47.765 153.810 ;
			LAYER M4 ;
			RECT 0.000 156.600 47.765 157.650 ;
			LAYER M4 ;
			RECT 0.000 160.440 47.765 160.940 ;
			LAYER M4 ;
			RECT 0.000 165.220 47.765 165.720 ;
			LAYER M4 ;
			RECT 0.000 167.110 47.765 167.610 ;
			LAYER M4 ;
			RECT 0.000 168.920 47.765 169.420 ;
			LAYER M4 ;
			RECT 0.000 169.550 47.765 169.950 ;
			LAYER M4 ;
			RECT 0.000 173.560 47.765 173.770 ;
			LAYER M4 ;
			RECT 32.420 173.870 47.765 174.110 ;
			LAYER M4 ;
			RECT 0.000 175.760 47.765 175.970 ;
			LAYER M4 ;
			RECT 32.420 176.070 47.765 176.310 ;
			LAYER M4 ;
			RECT 0.000 177.960 47.765 178.170 ;
			LAYER M4 ;
			RECT 32.420 178.270 47.765 178.490 ;
			LAYER M4 ;
			RECT 0.000 180.160 47.765 180.370 ;
			LAYER M4 ;
			RECT 32.420 180.470 47.765 180.710 ;
			LAYER M4 ;
			RECT 0.000 182.360 47.765 182.570 ;
			LAYER M4 ;
			RECT 32.420 182.670 47.765 182.890 ;
			LAYER M4 ;
			RECT 0.000 184.560 47.765 184.770 ;
			LAYER M4 ;
			RECT 32.420 184.870 47.765 185.110 ;
			LAYER M4 ;
			RECT 0.000 186.760 47.765 186.970 ;
			LAYER M4 ;
			RECT 32.420 187.070 47.765 187.290 ;
			LAYER M4 ;
			RECT 0.000 188.960 47.765 189.170 ;
			LAYER M4 ;
			RECT 32.420 189.270 47.765 189.510 ;
			LAYER M4 ;
			RECT 0.000 191.160 47.765 191.370 ;
			LAYER M4 ;
			RECT 32.420 191.470 47.765 191.690 ;
			LAYER M4 ;
			RECT 0.000 193.360 47.765 193.570 ;
			LAYER M4 ;
			RECT 32.420 193.670 47.765 193.910 ;
			LAYER M4 ;
			RECT 0.000 195.560 47.765 195.770 ;
			LAYER M4 ;
			RECT 32.420 195.870 47.765 196.090 ;
			LAYER M4 ;
			RECT 0.000 197.760 47.765 197.970 ;
			LAYER M4 ;
			RECT 32.420 198.070 47.765 198.310 ;
			LAYER M4 ;
			RECT 0.000 199.960 47.765 200.170 ;
			LAYER M4 ;
			RECT 32.420 200.270 47.765 200.490 ;
			LAYER M4 ;
			RECT 0.000 202.160 47.765 202.370 ;
			LAYER M4 ;
			RECT 32.420 202.470 47.765 202.710 ;
			LAYER M4 ;
			RECT 0.000 204.360 47.765 204.570 ;
			LAYER M4 ;
			RECT 32.420 204.670 47.765 204.890 ;
			LAYER M4 ;
			RECT 0.000 206.560 47.765 206.770 ;
			LAYER M4 ;
			RECT 32.420 206.870 47.765 207.110 ;
			LAYER M4 ;
			RECT 0.000 208.760 47.765 208.970 ;
			LAYER M4 ;
			RECT 32.420 209.070 47.765 209.290 ;
			LAYER M4 ;
			RECT 0.000 210.960 47.765 211.170 ;
			LAYER M4 ;
			RECT 32.420 211.270 47.765 211.510 ;
			LAYER M4 ;
			RECT 0.000 213.160 47.765 213.370 ;
			LAYER M4 ;
			RECT 32.420 213.470 47.765 213.690 ;
			LAYER M4 ;
			RECT 0.000 215.360 47.765 215.570 ;
			LAYER M4 ;
			RECT 32.420 215.670 47.765 215.910 ;
			LAYER M4 ;
			RECT 0.000 217.560 47.765 217.770 ;
			LAYER M4 ;
			RECT 32.420 217.870 47.765 218.090 ;
			LAYER M4 ;
			RECT 0.000 219.760 47.765 219.970 ;
			LAYER M4 ;
			RECT 32.420 220.070 47.765 220.310 ;
			LAYER M4 ;
			RECT 0.000 221.960 47.765 222.170 ;
			LAYER M4 ;
			RECT 32.420 222.270 47.765 222.490 ;
			LAYER M4 ;
			RECT 0.000 224.160 47.765 224.370 ;
			LAYER M4 ;
			RECT 32.420 224.470 47.765 224.710 ;
			LAYER M4 ;
			RECT 0.000 226.360 47.765 226.570 ;
			LAYER M4 ;
			RECT 32.420 226.670 47.765 226.890 ;
			LAYER M4 ;
			RECT 0.000 228.560 47.765 228.770 ;
			LAYER M4 ;
			RECT 32.420 228.870 47.765 229.110 ;
			LAYER M4 ;
			RECT 0.000 230.760 47.765 230.970 ;
			LAYER M4 ;
			RECT 32.420 231.070 47.765 231.290 ;
			LAYER M4 ;
			RECT 0.000 232.960 47.765 233.170 ;
			LAYER M4 ;
			RECT 32.420 233.270 47.765 233.510 ;
			LAYER M4 ;
			RECT 0.000 235.160 47.765 235.370 ;
			LAYER M4 ;
			RECT 32.420 235.470 47.765 235.690 ;
			LAYER M4 ;
			RECT 0.000 237.360 47.765 237.570 ;
			LAYER M4 ;
			RECT 32.420 237.670 47.765 237.910 ;
			LAYER M4 ;
			RECT 0.000 239.560 47.765 239.770 ;
			LAYER M4 ;
			RECT 32.420 239.870 47.765 240.090 ;
			LAYER M4 ;
			RECT 0.000 241.760 47.765 241.970 ;
			LAYER M4 ;
			RECT 32.420 242.070 47.765 242.310 ;
			LAYER M4 ;
			RECT 0.000 243.960 47.765 244.170 ;
			LAYER M4 ;
			RECT 32.420 244.270 47.765 244.490 ;
			LAYER M4 ;
			RECT 0.000 246.160 47.765 246.370 ;
			LAYER M4 ;
			RECT 32.420 246.470 47.765 246.710 ;
			LAYER M4 ;
			RECT 0.000 248.360 47.765 248.570 ;
			LAYER M4 ;
			RECT 32.420 248.670 47.765 248.890 ;
			LAYER M4 ;
			RECT 0.000 250.560 47.765 250.770 ;
			LAYER M4 ;
			RECT 32.420 250.870 47.765 251.110 ;
			LAYER M4 ;
			RECT 0.000 252.760 47.765 252.970 ;
			LAYER M4 ;
			RECT 32.420 253.070 47.765 253.290 ;
			LAYER M4 ;
			RECT 0.000 254.960 47.765 255.170 ;
			LAYER M4 ;
			RECT 32.420 255.270 47.765 255.510 ;
			LAYER M4 ;
			RECT 0.000 257.160 47.765 257.370 ;
			LAYER M4 ;
			RECT 32.420 257.470 47.765 257.690 ;
			LAYER M4 ;
			RECT 0.000 259.360 47.765 259.570 ;
			LAYER M4 ;
			RECT 32.420 259.670 47.765 259.910 ;
			LAYER M4 ;
			RECT 0.000 261.560 47.765 261.770 ;
			LAYER M4 ;
			RECT 32.420 261.870 47.765 262.090 ;
			LAYER M4 ;
			RECT 0.000 263.760 47.765 263.970 ;
			LAYER M4 ;
			RECT 32.420 264.070 47.765 264.310 ;
			LAYER M4 ;
			RECT 0.000 265.960 47.765 266.170 ;
			LAYER M4 ;
			RECT 32.420 266.270 47.765 266.490 ;
			LAYER M4 ;
			RECT 0.000 268.160 47.765 268.370 ;
			LAYER M4 ;
			RECT 32.420 268.470 47.765 268.710 ;
			LAYER M4 ;
			RECT 0.000 270.360 47.765 270.570 ;
			LAYER M4 ;
			RECT 32.420 270.670 47.765 270.890 ;
			LAYER M4 ;
			RECT 0.000 272.560 47.765 272.770 ;
			LAYER M4 ;
			RECT 32.420 272.870 47.765 273.110 ;
			LAYER M4 ;
			RECT 0.000 274.760 47.765 274.970 ;
			LAYER M4 ;
			RECT 32.420 275.070 47.765 275.290 ;
			LAYER M4 ;
			RECT 0.000 276.960 47.765 277.170 ;
			LAYER M4 ;
			RECT 32.420 277.270 47.765 277.510 ;
			LAYER M4 ;
			RECT 0.000 279.160 47.765 279.370 ;
			LAYER M4 ;
			RECT 32.420 279.470 47.765 279.690 ;
			LAYER M4 ;
			RECT 0.000 281.360 47.765 281.570 ;
			LAYER M4 ;
			RECT 32.420 281.670 47.765 281.910 ;
			LAYER M4 ;
			RECT 0.000 283.560 47.765 283.770 ;
			LAYER M4 ;
			RECT 32.420 283.870 47.765 284.090 ;
			LAYER M4 ;
			RECT 0.000 285.760 47.765 285.970 ;
			LAYER M4 ;
			RECT 32.420 286.070 47.765 286.310 ;
			LAYER M4 ;
			RECT 0.000 287.960 47.765 288.170 ;
			LAYER M4 ;
			RECT 32.420 288.270 47.765 288.490 ;
			LAYER M4 ;
			RECT 0.000 290.160 47.765 290.370 ;
			LAYER M4 ;
			RECT 32.420 290.470 47.765 290.710 ;
			LAYER M4 ;
			RECT 0.000 292.360 47.765 292.570 ;
			LAYER M4 ;
			RECT 32.420 292.670 47.765 292.890 ;
			LAYER M4 ;
			RECT 0.000 294.560 47.765 294.770 ;
			LAYER M4 ;
			RECT 32.420 294.870 47.765 295.110 ;
			LAYER M4 ;
			RECT 0.000 296.760 47.765 296.970 ;
			LAYER M4 ;
			RECT 32.420 297.070 47.765 297.290 ;
			LAYER M4 ;
			RECT 0.000 298.960 47.765 299.170 ;
			LAYER M4 ;
			RECT 32.420 299.270 47.765 299.510 ;
			LAYER M4 ;
			RECT 0.000 301.160 47.765 301.370 ;
			LAYER M4 ;
			RECT 32.420 301.470 47.765 301.690 ;
			LAYER M4 ;
			RECT 0.000 303.360 47.765 303.570 ;
			LAYER M4 ;
			RECT 32.420 303.670 47.765 303.910 ;
			LAYER M4 ;
			RECT 0.000 305.560 47.765 305.770 ;
			LAYER M4 ;
			RECT 32.420 305.870 47.765 306.090 ;
			LAYER M4 ;
			RECT 0.000 307.760 47.765 307.970 ;
			LAYER M4 ;
			RECT 32.420 308.070 47.765 308.310 ;
			LAYER M4 ;
			RECT 0.000 309.960 47.765 310.170 ;
			LAYER M4 ;
			RECT 32.420 310.270 47.765 310.490 ;
			LAYER M4 ;
			RECT 0.000 312.160 47.765 312.370 ;
			LAYER M4 ;
			RECT 32.420 312.470 47.765 312.710 ;
			LAYER M4 ;
			RECT 0.000 314.360 47.765 314.570 ;
			LAYER M4 ;
			RECT 32.420 314.670 47.765 314.890 ;
			LAYER M4 ;
			RECT 0.000 316.560 47.765 316.770 ;
		END
	END VSS

	PIN WCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 167.310 47.765 167.460 ;
			LAYER M2 ;
			RECT 47.525 167.310 47.765 167.460 ;
			LAYER M1 ;
			RECT 47.525 167.310 47.765 167.460 ;
		END
		ANTENNAGATEAREA 0.0308 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.2296 LAYER M1 ;
		ANTENNAMAXAREACAR 2.7922 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0280 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.3247 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0308 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.8892 LAYER M2 ;
		ANTENNAMAXAREACAR 30.8831 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0140 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.6981 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0308 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.1554 LAYER M3 ;
		ANTENNAMAXAREACAR 33.1315 LAYER M3 ;
	END WCT[0]

	PIN WCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.525 167.620 47.765 167.770 ;
			LAYER M3 ;
			RECT 47.525 167.620 47.765 167.770 ;
			LAYER M1 ;
			RECT 47.525 167.620 47.765 167.770 ;
		END
		ANTENNAGATEAREA 0.0308 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.2296 LAYER M1 ;
		ANTENNAMAXAREACAR 2.7922 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0280 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.3247 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0308 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.8892 LAYER M2 ;
		ANTENNAMAXAREACAR 30.8831 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0140 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.6981 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0308 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.1554 LAYER M3 ;
		ANTENNAMAXAREACAR 33.1315 LAYER M3 ;
	END WCT[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.525 163.610 47.765 163.760 ;
			LAYER M1 ;
			RECT 47.525 163.610 47.765 163.760 ;
			LAYER M2 ;
			RECT 47.525 163.610 47.765 163.760 ;
		END
		ANTENNAGATEAREA 0.0350 LAYER M1 ;
		ANTENNADIFFAREA 0.0350 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1953 LAYER M1 ;
		ANTENNAMAXAREACAR 4.5514 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0130 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.1857 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0350 LAYER M2 ;
		ANTENNADIFFAREA 0.0350 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0894 LAYER M2 ;
		ANTENNAMAXAREACAR 7.1057 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.3714 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0350 LAYER M3 ;
		ANTENNADIFFAREA 0.0350 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.0360 LAYER M3 ;
		ANTENNAMAXAREACAR 8.1343 LAYER M3 ;
	END WEB

	OBS
		# Promoted blockages
		LAYER M1 ;
		RECT 47.615 315.470 47.765 316.190 ;
		LAYER M3 ;
		RECT 47.615 312.230 47.765 315.030 ;
		LAYER M2 ;
		RECT 47.615 311.070 47.765 311.790 ;
		LAYER M3 ;
		RECT 47.615 311.070 47.765 311.790 ;
		LAYER M2 ;
		RECT 47.615 312.230 47.765 315.030 ;
		LAYER M2 ;
		RECT 47.615 315.470 47.765 316.190 ;
		LAYER M3 ;
		RECT 47.615 315.470 47.765 316.190 ;
		LAYER M1 ;
		RECT 47.615 311.070 47.765 311.790 ;
		LAYER M1 ;
		RECT 47.615 306.670 47.765 307.390 ;
		LAYER M1 ;
		RECT 47.615 303.430 47.765 306.230 ;
		LAYER M2 ;
		RECT 47.615 303.430 47.765 306.230 ;
		LAYER M3 ;
		RECT 47.615 307.830 47.765 310.630 ;
		LAYER M3 ;
		RECT 47.615 303.430 47.765 306.230 ;
		LAYER M2 ;
		RECT 47.615 306.670 47.765 307.390 ;
		LAYER M3 ;
		RECT 47.615 306.670 47.765 307.390 ;
		LAYER M2 ;
		RECT 47.615 307.830 47.765 310.630 ;
		LAYER M1 ;
		RECT 47.615 307.830 47.765 310.630 ;
		LAYER M1 ;
		RECT 47.615 297.870 47.765 298.590 ;
		LAYER M1 ;
		RECT 47.615 299.030 47.765 301.830 ;
		LAYER M2 ;
		RECT 47.615 299.030 47.765 301.830 ;
		LAYER M3 ;
		RECT 47.615 299.030 47.765 301.830 ;
		LAYER M2 ;
		RECT 47.615 297.870 47.765 298.590 ;
		LAYER M3 ;
		RECT 47.615 297.870 47.765 298.590 ;
		LAYER M1 ;
		RECT 47.615 302.270 47.765 302.990 ;
		LAYER M2 ;
		RECT 47.615 302.270 47.765 302.990 ;
		LAYER M3 ;
		RECT 47.615 302.270 47.765 302.990 ;
		LAYER M1 ;
		RECT 47.615 294.630 47.765 297.430 ;
		LAYER M3 ;
		RECT 47.615 290.230 47.765 293.030 ;
		LAYER M1 ;
		RECT 47.615 290.230 47.765 293.030 ;
		LAYER M2 ;
		RECT 47.615 294.630 47.765 297.430 ;
		LAYER M3 ;
		RECT 47.615 294.630 47.765 297.430 ;
		LAYER M1 ;
		RECT 47.615 289.070 47.765 289.790 ;
		LAYER M2 ;
		RECT 47.615 289.070 47.765 289.790 ;
		LAYER M3 ;
		RECT 47.615 289.070 47.765 289.790 ;
		LAYER M2 ;
		RECT 47.615 293.470 47.765 294.190 ;
		LAYER M3 ;
		RECT 47.615 293.470 47.765 294.190 ;
		LAYER M1 ;
		RECT 47.615 293.470 47.765 294.190 ;
		LAYER M2 ;
		RECT 47.615 290.230 47.765 293.030 ;
		LAYER M1 ;
		RECT 47.615 285.830 47.765 288.630 ;
		LAYER M2 ;
		RECT 47.615 284.670 47.765 285.390 ;
		LAYER M3 ;
		RECT 47.615 284.670 47.765 285.390 ;
		LAYER M2 ;
		RECT 47.615 281.430 47.765 284.230 ;
		LAYER M1 ;
		RECT 47.615 284.670 47.765 285.390 ;
		LAYER M1 ;
		RECT 47.615 281.430 47.765 284.230 ;
		LAYER M3 ;
		RECT 47.615 277.030 47.765 279.830 ;
		LAYER M3 ;
		RECT 47.615 275.870 47.765 276.590 ;
		LAYER M2 ;
		RECT 47.615 275.870 47.765 276.590 ;
		LAYER M1 ;
		RECT 47.615 280.270 47.765 280.990 ;
		LAYER M1 ;
		RECT 47.615 275.870 47.765 276.590 ;
		LAYER M3 ;
		RECT 47.615 271.470 47.765 272.190 ;
		LAYER M3 ;
		RECT 47.615 272.630 47.765 275.430 ;
		LAYER M1 ;
		RECT 47.615 272.630 47.765 275.430 ;
		LAYER M1 ;
		RECT 47.615 268.230 47.765 271.030 ;
		LAYER M2 ;
		RECT 47.615 272.630 47.765 275.430 ;
		LAYER M2 ;
		RECT 47.615 285.830 47.765 288.630 ;
		LAYER M3 ;
		RECT 47.615 285.830 47.765 288.630 ;
		LAYER M3 ;
		RECT 47.615 281.430 47.765 284.230 ;
		LAYER M1 ;
		RECT 47.615 277.030 47.765 279.830 ;
		LAYER M2 ;
		RECT 47.615 277.030 47.765 279.830 ;
		LAYER M2 ;
		RECT 47.615 280.270 47.765 280.990 ;
		LAYER M3 ;
		RECT 47.615 280.270 47.765 280.990 ;
		LAYER M1 ;
		RECT 47.615 271.470 47.765 272.190 ;
		LAYER M1 ;
		RECT 47.615 267.070 47.765 267.790 ;
		LAYER M3 ;
		RECT 47.615 267.070 47.765 267.790 ;
		LAYER M2 ;
		RECT 47.615 271.470 47.765 272.190 ;
		LAYER M3 ;
		RECT 47.615 268.230 47.765 271.030 ;
		LAYER M1 ;
		RECT 47.615 253.870 47.765 254.590 ;
		LAYER M2 ;
		RECT 47.615 255.030 47.765 257.830 ;
		LAYER M3 ;
		RECT 47.615 255.030 47.765 257.830 ;
		LAYER M1 ;
		RECT 47.615 258.270 47.765 258.990 ;
		LAYER M1 ;
		RECT 47.615 255.030 47.765 257.830 ;
		LAYER M3 ;
		RECT 47.615 253.870 47.765 254.590 ;
		LAYER M1 ;
		RECT 47.615 249.470 47.765 250.190 ;
		LAYER M2 ;
		RECT 47.615 249.470 47.765 250.190 ;
		LAYER M1 ;
		RECT 47.615 250.630 47.765 253.430 ;
		LAYER M2 ;
		RECT 47.615 250.630 47.765 253.430 ;
		LAYER M3 ;
		RECT 47.615 250.630 47.765 253.430 ;
		LAYER M3 ;
		RECT 47.615 249.470 47.765 250.190 ;
		LAYER M3 ;
		RECT 47.615 246.230 47.765 249.030 ;
		LAYER M1 ;
		RECT 47.615 246.230 47.765 249.030 ;
		LAYER M2 ;
		RECT 47.615 246.230 47.765 249.030 ;
		LAYER M1 ;
		RECT 47.615 245.070 47.765 245.790 ;
		LAYER M1 ;
		RECT 47.615 263.830 47.765 266.630 ;
		LAYER M3 ;
		RECT 47.615 263.830 47.765 266.630 ;
		LAYER M2 ;
		RECT 47.615 263.830 47.765 266.630 ;
		LAYER M2 ;
		RECT 47.615 253.870 47.765 254.590 ;
		LAYER M2 ;
		RECT 47.615 258.270 47.765 258.990 ;
		LAYER M3 ;
		RECT 47.615 258.270 47.765 258.990 ;
		LAYER M1 ;
		RECT 47.615 259.430 47.765 262.230 ;
		LAYER M2 ;
		RECT 47.615 259.430 47.765 262.230 ;
		LAYER M3 ;
		RECT 47.615 259.430 47.765 262.230 ;
		LAYER M1 ;
		RECT 47.615 262.670 47.765 263.390 ;
		LAYER M3 ;
		RECT 47.615 262.670 47.765 263.390 ;
		LAYER M2 ;
		RECT 47.615 262.670 47.765 263.390 ;
		LAYER M1 ;
		RECT 47.615 21.655 47.765 22.375 ;
		LAYER M3 ;
		RECT 47.615 21.655 47.765 22.375 ;
		LAYER M2 ;
		RECT 47.615 49.215 47.765 52.015 ;
		LAYER M1 ;
		RECT 47.615 31.615 47.765 34.415 ;
		LAYER M1 ;
		RECT 47.615 43.655 47.765 44.375 ;
		LAYER M3 ;
		RECT 47.615 44.815 47.765 47.615 ;
		LAYER M2 ;
		RECT 47.615 61.255 47.765 61.975 ;
		LAYER M1 ;
		RECT 47.615 58.015 47.765 60.815 ;
		LAYER M2 ;
		RECT 47.615 62.415 47.765 65.215 ;
		LAYER M3 ;
		RECT 47.615 62.415 47.765 65.215 ;
		LAYER M3 ;
		RECT 47.615 61.255 47.765 61.975 ;
		LAYER M1 ;
		RECT 47.615 61.255 47.765 61.975 ;
		LAYER M1 ;
		RECT 47.615 40.415 47.765 43.215 ;
		LAYER M2 ;
		RECT 47.615 40.415 47.765 43.215 ;
		LAYER M3 ;
		RECT 47.615 40.415 47.765 43.215 ;
		LAYER M2 ;
		RECT 47.615 65.655 47.765 66.375 ;
		LAYER M3 ;
		RECT 47.615 65.655 47.765 66.375 ;
		LAYER M3 ;
		RECT 47.615 66.815 47.765 69.615 ;
		LAYER M3 ;
		RECT 47.615 56.855 47.765 57.575 ;
		LAYER M3 ;
		RECT 47.615 70.055 47.765 70.775 ;
		LAYER M2 ;
		RECT 47.615 52.455 47.765 53.175 ;
		LAYER M3 ;
		RECT 47.615 52.455 47.765 53.175 ;
		LAYER M2 ;
		RECT 47.615 53.615 47.765 56.415 ;
		LAYER M3 ;
		RECT 47.615 53.615 47.765 56.415 ;
		LAYER M1 ;
		RECT 47.615 22.815 47.765 25.615 ;
		LAYER M2 ;
		RECT 47.615 22.815 47.765 25.615 ;
		LAYER M3 ;
		RECT 47.615 22.815 47.765 25.615 ;
		LAYER M1 ;
		RECT 47.615 48.055 47.765 48.775 ;
		LAYER M1 ;
		RECT 47.615 44.815 47.765 47.615 ;
		LAYER M2 ;
		RECT 47.615 44.815 47.765 47.615 ;
		LAYER M2 ;
		RECT 47.615 43.655 47.765 44.375 ;
		LAYER M2 ;
		RECT 47.615 39.255 47.765 39.975 ;
		LAYER M3 ;
		RECT 47.615 39.255 47.765 39.975 ;
		LAYER M2 ;
		RECT 47.615 36.015 47.765 38.815 ;
		LAYER M3 ;
		RECT 47.615 36.015 47.765 38.815 ;
		LAYER M3 ;
		RECT 47.615 34.855 47.765 35.575 ;
		LAYER M1 ;
		RECT 47.615 26.055 47.765 26.775 ;
		LAYER M2 ;
		RECT 47.615 26.055 47.765 26.775 ;
		LAYER M3 ;
		RECT 47.615 26.055 47.765 26.775 ;
		LAYER M1 ;
		RECT 47.615 27.215 47.765 30.015 ;
		LAYER M3 ;
		RECT 47.615 27.215 47.765 30.015 ;
		LAYER M2 ;
		RECT 47.615 27.215 47.765 30.015 ;
		LAYER M3 ;
		RECT 47.615 30.455 47.765 31.175 ;
		LAYER M2 ;
		RECT 47.615 48.055 47.765 48.775 ;
		LAYER M3 ;
		RECT 47.615 48.055 47.765 48.775 ;
		LAYER M3 ;
		RECT 47.615 43.655 47.765 44.375 ;
		LAYER M1 ;
		RECT 47.615 87.655 47.765 88.375 ;
		LAYER M2 ;
		RECT 47.615 84.415 47.765 87.215 ;
		LAYER M3 ;
		RECT 47.615 84.415 47.765 87.215 ;
		LAYER M2 ;
		RECT 47.615 87.655 47.765 88.375 ;
		LAYER M3 ;
		RECT 47.615 87.655 47.765 88.375 ;
		LAYER M1 ;
		RECT 47.615 84.415 47.765 87.215 ;
		LAYER M1 ;
		RECT 47.615 83.255 47.765 83.975 ;
		LAYER M2 ;
		RECT 47.615 78.855 47.765 79.575 ;
		LAYER M3 ;
		RECT 47.615 78.855 47.765 79.575 ;
		LAYER M2 ;
		RECT 47.615 83.255 47.765 83.975 ;
		LAYER M3 ;
		RECT 47.615 75.615 47.765 78.415 ;
		LAYER M1 ;
		RECT 47.615 75.615 47.765 78.415 ;
		LAYER M2 ;
		RECT 47.615 75.615 47.765 78.415 ;
		LAYER M1 ;
		RECT 47.615 80.015 47.765 82.815 ;
		LAYER M2 ;
		RECT 47.615 80.015 47.765 82.815 ;
		LAYER M3 ;
		RECT 47.615 80.015 47.765 82.815 ;
		LAYER M1 ;
		RECT 47.615 78.855 47.765 79.575 ;
		LAYER M3 ;
		RECT 47.615 83.255 47.765 83.975 ;
		LAYER M3 ;
		RECT 47.615 74.455 47.765 75.175 ;
		LAYER M3 ;
		RECT 47.615 71.215 47.765 74.015 ;
		LAYER M1 ;
		RECT 47.615 88.815 47.765 91.615 ;
		LAYER M2 ;
		RECT 47.615 97.615 47.765 100.415 ;
		LAYER M3 ;
		RECT 47.615 97.615 47.765 100.415 ;
		LAYER M3 ;
		RECT 47.615 88.815 47.765 91.615 ;
		LAYER M2 ;
		RECT 47.615 88.815 47.765 91.615 ;
		LAYER M3 ;
		RECT 47.615 96.455 47.765 97.175 ;
		LAYER M2 ;
		RECT 47.615 92.055 47.765 92.775 ;
		LAYER M2 ;
		RECT 47.615 93.215 47.765 96.015 ;
		LAYER M3 ;
		RECT 47.615 93.215 47.765 96.015 ;
		LAYER M2 ;
		RECT 47.615 96.455 47.765 97.175 ;
		LAYER M2 ;
		RECT 47.615 105.255 47.765 105.975 ;
		LAYER M3 ;
		RECT 47.615 105.255 47.765 105.975 ;
		LAYER M1 ;
		RECT 47.615 105.255 47.765 105.975 ;
		LAYER M3 ;
		RECT 47.615 106.415 47.765 109.215 ;
		LAYER M2 ;
		RECT 47.615 106.415 47.765 109.215 ;
		LAYER M1 ;
		RECT 47.615 312.230 47.765 315.030 ;
		LAYER M1 ;
		RECT 47.615 36.015 47.765 38.815 ;
		LAYER M1 ;
		RECT 47.615 4.055 47.765 4.775 ;
		LAYER M1 ;
		RECT 47.615 65.655 47.765 66.375 ;
		LAYER M1 ;
		RECT 47.615 62.415 47.765 65.215 ;
		LAYER M1 ;
		RECT 47.615 39.255 47.765 39.975 ;
		LAYER M1 ;
		RECT 47.615 316.630 47.765 317.515 ;
		LAYER M2 ;
		RECT 47.615 316.630 47.765 317.515 ;
		LAYER M3 ;
		RECT 47.615 316.630 47.765 317.515 ;
		LAYER M1 ;
		RECT 47.525 173.400 47.615 317.515 ;
		LAYER M2 ;
		RECT 47.525 173.420 47.615 317.515 ;
		LAYER M3 ;
		RECT 47.525 146.915 47.765 149.245 ;
		LAYER M1 ;
		RECT 47.525 146.585 47.765 146.625 ;
		LAYER M3 ;
		RECT 47.525 173.420 47.615 317.515 ;
		LAYER M1 ;
		RECT 47.525 0.000 47.615 146.315 ;
		LAYER M3 ;
		RECT 47.525 0.000 47.615 146.295 ;
		LAYER M2 ;
		RECT 47.525 0.000 47.615 146.295 ;
		LAYER M1 ;
		RECT 0.000 0.000 47.525 317.515 ;
		LAYER M2 ;
		RECT 0.000 0.000 47.525 317.515 ;
		LAYER M3 ;
		RECT 0.000 0.000 47.525 317.515 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 47.765 317.515 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 47.765 317.515 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 47.765 317.515 ;
		LAYER M2 ;
		RECT 47.615 21.655 47.765 22.375 ;
		LAYER M2 ;
		RECT 47.615 31.615 47.765 34.415 ;
		LAYER M3 ;
		RECT 47.615 31.615 47.765 34.415 ;
		LAYER M2 ;
		RECT 47.615 34.855 47.765 35.575 ;
		LAYER M1 ;
		RECT 47.615 34.855 47.765 35.575 ;
		LAYER M1 ;
		RECT 47.615 30.455 47.765 31.175 ;
		LAYER M2 ;
		RECT 47.615 30.455 47.765 31.175 ;
		LAYER M2 ;
		RECT 47.615 18.415 47.765 21.215 ;
		LAYER M3 ;
		RECT 47.615 18.415 47.765 21.215 ;
		LAYER M1 ;
		RECT 47.615 56.855 47.765 57.575 ;
		LAYER M2 ;
		RECT 47.615 56.855 47.765 57.575 ;
		LAYER M1 ;
		RECT 47.615 53.615 47.765 56.415 ;
		LAYER M1 ;
		RECT 47.615 52.455 47.765 53.175 ;
		LAYER M2 ;
		RECT 47.615 66.815 47.765 69.615 ;
		LAYER M1 ;
		RECT 47.615 49.215 47.765 52.015 ;
		LAYER M3 ;
		RECT 47.615 49.215 47.765 52.015 ;
		LAYER M2 ;
		RECT 47.615 4.055 47.765 4.775 ;
		LAYER M3 ;
		RECT 47.615 4.055 47.765 4.775 ;
		LAYER M2 ;
		RECT 47.615 5.215 47.765 8.015 ;
		LAYER M1 ;
		RECT 47.615 5.215 47.765 8.015 ;
		LAYER M3 ;
		RECT 47.615 5.215 47.765 8.015 ;
		LAYER M1 ;
		RECT 47.615 106.415 47.765 109.215 ;
		LAYER M3 ;
		RECT 47.615 102.015 47.765 104.815 ;
		LAYER M1 ;
		RECT 47.615 102.015 47.765 104.815 ;
		LAYER M3 ;
		RECT 47.615 245.070 47.765 245.790 ;
		LAYER M3 ;
		RECT 47.615 237.430 47.765 240.230 ;
		LAYER M1 ;
		RECT 47.615 8.455 47.765 9.175 ;
		LAYER M1 ;
		RECT 47.615 140.455 47.765 141.175 ;
		LAYER M1 ;
		RECT 47.615 127.255 47.765 127.975 ;
		LAYER M2 ;
		RECT 47.615 127.255 47.765 127.975 ;
		LAYER M1 ;
		RECT 47.525 158.230 47.765 161.950 ;
		LAYER M2 ;
		RECT 47.525 158.250 47.765 161.930 ;
		LAYER M1 ;
		RECT 47.525 157.920 47.765 157.960 ;
		LAYER M2 ;
		RECT 47.525 157.320 47.765 157.630 ;
		LAYER M1 ;
		RECT 47.525 156.165 47.765 157.030 ;
		LAYER M2 ;
		RECT 47.525 155.565 47.765 155.875 ;
		LAYER M3 ;
		RECT 47.525 155.565 47.765 155.875 ;
		LAYER M1 ;
		RECT 47.615 14.015 47.765 16.815 ;
		LAYER M1 ;
		RECT 47.615 17.255 47.765 17.975 ;
		LAYER M2 ;
		RECT 47.615 17.255 47.765 17.975 ;
		LAYER M3 ;
		RECT 47.615 17.255 47.765 17.975 ;
		LAYER M1 ;
		RECT 47.615 66.815 47.765 69.615 ;
		LAYER M1 ;
		RECT 47.615 70.055 47.765 70.775 ;
		LAYER M2 ;
		RECT 47.615 70.055 47.765 70.775 ;
		LAYER M2 ;
		RECT 47.615 58.015 47.765 60.815 ;
		LAYER M3 ;
		RECT 47.615 58.015 47.765 60.815 ;
		LAYER M1 ;
		RECT 47.615 74.455 47.765 75.175 ;
		LAYER M2 ;
		RECT 47.615 74.455 47.765 75.175 ;
		LAYER M1 ;
		RECT 47.615 71.215 47.765 74.015 ;
		LAYER M2 ;
		RECT 47.615 71.215 47.765 74.015 ;
		LAYER M2 ;
		RECT 47.615 14.015 47.765 16.815 ;
		LAYER M3 ;
		RECT 47.615 14.015 47.765 16.815 ;
		LAYER M1 ;
		RECT 47.615 18.415 47.765 21.215 ;
		LAYER M1 ;
		RECT 47.615 0.000 47.765 3.615 ;
		LAYER M2 ;
		RECT 47.615 0.000 47.765 3.615 ;
		LAYER M3 ;
		RECT 47.615 0.000 47.765 3.615 ;
		LAYER M3 ;
		RECT 47.615 8.455 47.765 9.175 ;
		LAYER M2 ;
		RECT 47.615 8.455 47.765 9.175 ;
		LAYER M1 ;
		RECT 47.615 9.615 47.765 12.415 ;
		LAYER M2 ;
		RECT 47.615 9.615 47.765 12.415 ;
		LAYER M1 ;
		RECT 47.615 12.855 47.765 13.575 ;
		LAYER M3 ;
		RECT 47.615 12.855 47.765 13.575 ;
		LAYER M3 ;
		RECT 47.615 9.615 47.765 12.415 ;
		LAYER M1 ;
		RECT 47.615 92.055 47.765 92.775 ;
		LAYER M2 ;
		RECT 47.615 12.855 47.765 13.575 ;
		LAYER M1 ;
		RECT 47.615 97.615 47.765 100.415 ;
		LAYER M1 ;
		RECT 47.615 96.455 47.765 97.175 ;
		LAYER M1 ;
		RECT 47.615 93.215 47.765 96.015 ;
		LAYER M3 ;
		RECT 47.615 92.055 47.765 92.775 ;
		LAYER M2 ;
		RECT 47.615 100.855 47.765 101.575 ;
		LAYER M3 ;
		RECT 47.615 100.855 47.765 101.575 ;
		LAYER M1 ;
		RECT 47.615 100.855 47.765 101.575 ;
		LAYER M2 ;
		RECT 47.615 102.015 47.765 104.815 ;
		LAYER M1 ;
		RECT 47.615 228.630 47.765 231.430 ;
		LAYER M3 ;
		RECT 47.615 227.470 47.765 228.190 ;
		LAYER M1 ;
		RECT 47.615 227.470 47.765 228.190 ;
		LAYER M2 ;
		RECT 47.615 231.870 47.765 232.590 ;
		LAYER M2 ;
		RECT 47.615 183.470 47.765 184.190 ;
		LAYER M1 ;
		RECT 47.615 180.230 47.765 183.030 ;
		LAYER M1 ;
		RECT 47.615 179.070 47.765 179.790 ;
		LAYER M2 ;
		RECT 47.615 179.070 47.765 179.790 ;
		LAYER M2 ;
		RECT 47.615 180.230 47.765 183.030 ;
		LAYER M3 ;
		RECT 47.615 180.230 47.765 183.030 ;
		LAYER M3 ;
		RECT 47.615 179.070 47.765 179.790 ;
		LAYER M1 ;
		RECT 47.615 141.615 47.765 146.315 ;
		LAYER M2 ;
		RECT 47.615 141.615 47.765 146.295 ;
		LAYER M3 ;
		RECT 47.615 173.420 47.765 178.630 ;
		LAYER M1 ;
		RECT 47.615 173.400 47.765 178.630 ;
		LAYER M2 ;
		RECT 47.615 173.420 47.765 178.630 ;
		LAYER M3 ;
		RECT 47.615 206.630 47.765 209.430 ;
		LAYER M3 ;
		RECT 47.615 122.855 47.765 123.575 ;
		LAYER M3 ;
		RECT 47.615 118.455 47.765 119.175 ;
		LAYER M2 ;
		RECT 47.615 119.615 47.765 122.415 ;
		LAYER M1 ;
		RECT 47.615 119.615 47.765 122.415 ;
		LAYER M3 ;
		RECT 47.615 119.615 47.765 122.415 ;
		LAYER M1 ;
		RECT 47.615 115.215 47.765 118.015 ;
		LAYER M2 ;
		RECT 47.615 115.215 47.765 118.015 ;
		LAYER M1 ;
		RECT 47.615 118.455 47.765 119.175 ;
		LAYER M2 ;
		RECT 47.615 118.455 47.765 119.175 ;
		LAYER M3 ;
		RECT 47.615 115.215 47.765 118.015 ;
		LAYER M2 ;
		RECT 47.615 245.070 47.765 245.790 ;
		LAYER M1 ;
		RECT 47.615 241.830 47.765 244.630 ;
		LAYER M2 ;
		RECT 47.615 241.830 47.765 244.630 ;
		LAYER M3 ;
		RECT 47.615 241.830 47.765 244.630 ;
		LAYER M2 ;
		RECT 47.615 267.070 47.765 267.790 ;
		LAYER M1 ;
		RECT 47.615 240.670 47.765 241.390 ;
		LAYER M2 ;
		RECT 47.615 240.670 47.765 241.390 ;
		LAYER M3 ;
		RECT 47.615 240.670 47.765 241.390 ;
		LAYER M1 ;
		RECT 47.615 124.015 47.765 126.815 ;
		LAYER M2 ;
		RECT 47.615 124.015 47.765 126.815 ;
		LAYER M3 ;
		RECT 47.615 124.015 47.765 126.815 ;
		LAYER M1 ;
		RECT 47.615 122.855 47.765 123.575 ;
		LAYER M3 ;
		RECT 47.615 132.815 47.765 135.615 ;
		LAYER M2 ;
		RECT 47.615 136.055 47.765 136.775 ;
		LAYER M3 ;
		RECT 47.615 136.055 47.765 136.775 ;
		LAYER M2 ;
		RECT 47.615 137.215 47.765 140.015 ;
		LAYER M2 ;
		RECT 47.615 132.815 47.765 135.615 ;
		LAYER M1 ;
		RECT 47.615 132.815 47.765 135.615 ;
		LAYER M2 ;
		RECT 47.615 140.455 47.765 141.175 ;
		LAYER M3 ;
		RECT 47.615 137.215 47.765 140.015 ;
		LAYER M2 ;
		RECT 47.615 122.855 47.765 123.575 ;
		LAYER M3 ;
		RECT 47.615 127.255 47.765 127.975 ;
		LAYER M1 ;
		RECT 47.615 128.415 47.765 131.215 ;
		LAYER M1 ;
		RECT 47.615 131.655 47.765 132.375 ;
		LAYER M3 ;
		RECT 47.615 131.655 47.765 132.375 ;
		LAYER M3 ;
		RECT 47.615 141.615 47.765 146.295 ;
		LAYER M3 ;
		RECT 47.615 140.455 47.765 141.175 ;
		LAYER M2 ;
		RECT 47.615 131.655 47.765 132.375 ;
		LAYER M1 ;
		RECT 47.615 109.655 47.765 110.375 ;
		LAYER M2 ;
		RECT 47.615 110.815 47.765 113.615 ;
		LAYER M3 ;
		RECT 47.615 110.815 47.765 113.615 ;
		LAYER M1 ;
		RECT 47.615 110.815 47.765 113.615 ;
		LAYER M2 ;
		RECT 47.615 109.655 47.765 110.375 ;
		LAYER M3 ;
		RECT 47.615 109.655 47.765 110.375 ;
		LAYER M1 ;
		RECT 47.615 114.055 47.765 114.775 ;
		LAYER M2 ;
		RECT 47.615 114.055 47.765 114.775 ;
		LAYER M3 ;
		RECT 47.615 114.055 47.765 114.775 ;
		LAYER M2 ;
		RECT 47.615 268.230 47.765 271.030 ;
		LAYER M1 ;
		RECT 47.615 237.430 47.765 240.230 ;
		LAYER M2 ;
		RECT 47.615 237.430 47.765 240.230 ;
		LAYER M3 ;
		RECT 47.615 228.630 47.765 231.430 ;
		LAYER M1 ;
		RECT 47.615 233.030 47.765 235.830 ;
		LAYER M2 ;
		RECT 47.615 233.030 47.765 235.830 ;
		LAYER M1 ;
		RECT 47.615 231.870 47.765 232.590 ;
		LAYER M3 ;
		RECT 47.615 231.870 47.765 232.590 ;
		LAYER M2 ;
		RECT 47.615 192.270 47.765 192.990 ;
		LAYER M1 ;
		RECT 47.615 184.630 47.765 187.430 ;
		LAYER M2 ;
		RECT 47.615 184.630 47.765 187.430 ;
		LAYER M3 ;
		RECT 47.615 184.630 47.765 187.430 ;
		LAYER M1 ;
		RECT 47.615 201.070 47.765 201.790 ;
		LAYER M1 ;
		RECT 47.615 183.470 47.765 184.190 ;
		LAYER M3 ;
		RECT 47.615 183.470 47.765 184.190 ;
		LAYER M3 ;
		RECT 47.615 233.030 47.765 235.830 ;
		LAYER M3 ;
		RECT 47.615 209.870 47.765 210.590 ;
		LAYER M2 ;
		RECT 47.615 209.870 47.765 210.590 ;
		LAYER M1 ;
		RECT 47.615 218.670 47.765 219.390 ;
		LAYER M2 ;
		RECT 47.615 218.670 47.765 219.390 ;
		LAYER M3 ;
		RECT 47.615 215.430 47.765 218.230 ;
		LAYER M1 ;
		RECT 47.615 209.870 47.765 210.590 ;
		LAYER M1 ;
		RECT 47.615 189.030 47.765 191.830 ;
		LAYER M2 ;
		RECT 47.615 189.030 47.765 191.830 ;
		LAYER M1 ;
		RECT 47.615 187.870 47.765 188.590 ;
		LAYER M2 ;
		RECT 47.615 187.870 47.765 188.590 ;
		LAYER M3 ;
		RECT 47.615 189.030 47.765 191.830 ;
		LAYER M3 ;
		RECT 47.615 187.870 47.765 188.590 ;
		LAYER M1 ;
		RECT 47.615 202.230 47.765 205.030 ;
		LAYER M2 ;
		RECT 47.615 201.070 47.765 201.790 ;
		LAYER M3 ;
		RECT 47.615 201.070 47.765 201.790 ;
		LAYER M1 ;
		RECT 47.615 197.830 47.765 200.630 ;
		LAYER M2 ;
		RECT 47.615 202.230 47.765 205.030 ;
		LAYER M3 ;
		RECT 47.615 202.230 47.765 205.030 ;
		LAYER M1 ;
		RECT 47.615 196.670 47.765 197.390 ;
		LAYER M2 ;
		RECT 47.615 197.830 47.765 200.630 ;
		LAYER M3 ;
		RECT 47.615 196.670 47.765 197.390 ;
		LAYER M2 ;
		RECT 47.615 196.670 47.765 197.390 ;
		LAYER M1 ;
		RECT 47.615 192.270 47.765 192.990 ;
		LAYER M3 ;
		RECT 47.615 192.270 47.765 192.990 ;
		LAYER M1 ;
		RECT 47.615 193.430 47.765 196.230 ;
		LAYER M3 ;
		RECT 47.615 193.430 47.765 196.230 ;
		LAYER M2 ;
		RECT 47.615 193.430 47.765 196.230 ;
		LAYER M2 ;
		RECT 47.615 205.470 47.765 206.190 ;
		LAYER M1 ;
		RECT 47.615 205.470 47.765 206.190 ;
		LAYER M3 ;
		RECT 47.615 197.830 47.765 200.630 ;
		LAYER M3 ;
		RECT 47.615 205.470 47.765 206.190 ;
		LAYER M1 ;
		RECT 47.615 236.270 47.765 236.990 ;
		LAYER M1 ;
		RECT 47.615 224.230 47.765 227.030 ;
		LAYER M2 ;
		RECT 47.615 224.230 47.765 227.030 ;
		LAYER M3 ;
		RECT 47.615 224.230 47.765 227.030 ;
		LAYER M2 ;
		RECT 47.615 228.630 47.765 231.430 ;
		LAYER M2 ;
		RECT 47.615 227.470 47.765 228.190 ;
		LAYER M1 ;
		RECT 47.615 215.430 47.765 218.230 ;
		LAYER M1 ;
		RECT 47.615 219.830 47.765 222.630 ;
		LAYER M3 ;
		RECT 47.615 219.830 47.765 222.630 ;
		LAYER M1 ;
		RECT 47.615 223.070 47.765 223.790 ;
		LAYER M2 ;
		RECT 47.615 219.830 47.765 222.630 ;
		LAYER M3 ;
		RECT 47.615 218.670 47.765 219.390 ;
		LAYER M2 ;
		RECT 47.615 236.270 47.765 236.990 ;
		LAYER M3 ;
		RECT 47.615 236.270 47.765 236.990 ;
		LAYER M2 ;
		RECT 47.615 206.630 47.765 209.430 ;
		LAYER M1 ;
		RECT 47.615 206.630 47.765 209.430 ;
		LAYER M1 ;
		RECT 47.615 214.270 47.765 214.990 ;
		LAYER M2 ;
		RECT 47.615 214.270 47.765 214.990 ;
		LAYER M2 ;
		RECT 47.615 215.430 47.765 218.230 ;
		LAYER M3 ;
		RECT 47.615 223.070 47.765 223.790 ;
		LAYER M2 ;
		RECT 47.615 223.070 47.765 223.790 ;
		LAYER M3 ;
		RECT 47.615 211.030 47.765 213.830 ;
		LAYER M1 ;
		RECT 47.615 211.030 47.765 213.830 ;
		LAYER M2 ;
		RECT 47.615 211.030 47.765 213.830 ;
		LAYER M3 ;
		RECT 47.615 214.270 47.765 214.990 ;
		LAYER M1 ;
		RECT 47.615 137.215 47.765 140.015 ;
		LAYER M1 ;
		RECT 47.615 136.055 47.765 136.775 ;
		LAYER M2 ;
		RECT 47.615 128.415 47.765 131.215 ;
		LAYER M3 ;
		RECT 47.615 128.415 47.765 131.215 ;
		LAYER M1 ;
		RECT 47.525 155.545 47.765 155.895 ;
		LAYER M2 ;
		RECT 47.525 156.185 47.765 157.010 ;
		LAYER M2 ;
		RECT 47.525 162.240 47.765 163.530 ;
		LAYER M3 ;
		RECT 47.525 156.185 47.765 157.010 ;
		LAYER M1 ;
		RECT 47.525 154.365 47.765 155.275 ;
		LAYER M3 ;
		RECT 47.525 163.840 47.765 165.330 ;
		LAYER M1 ;
		RECT 47.525 162.220 47.765 163.550 ;
		LAYER M3 ;
		RECT 47.525 157.320 47.765 157.630 ;
		LAYER M1 ;
		RECT 47.525 157.300 47.765 157.650 ;
		LAYER M3 ;
		RECT 47.525 158.250 47.765 161.930 ;
		LAYER M3 ;
		RECT 47.525 162.240 47.765 163.530 ;
		LAYER M2 ;
		RECT 47.525 146.915 47.765 149.245 ;
		LAYER M1 ;
		RECT 47.525 146.895 47.765 149.265 ;
		LAYER M2 ;
		RECT 47.525 149.555 47.765 150.185 ;
		LAYER M1 ;
		RECT 47.525 149.535 47.765 150.205 ;
		LAYER M1 ;
		RECT 47.525 150.475 47.765 150.515 ;
		LAYER M3 ;
		RECT 47.525 149.555 47.765 150.185 ;
		LAYER M1 ;
		RECT 47.525 151.715 47.765 152.845 ;
		LAYER M1 ;
		RECT 47.525 153.115 47.765 153.155 ;
		LAYER M1 ;
		RECT 47.525 151.405 47.765 151.445 ;
		LAYER M2 ;
		RECT 47.525 153.445 47.765 154.075 ;
		LAYER M3 ;
		RECT 47.525 151.735 47.765 152.825 ;
		LAYER M2 ;
		RECT 47.525 151.735 47.765 152.825 ;
		LAYER M2 ;
		RECT 47.525 150.805 47.765 151.115 ;
		LAYER M1 ;
		RECT 47.525 153.425 47.765 154.095 ;
		LAYER M3 ;
		RECT 47.525 153.445 47.765 154.075 ;
		LAYER M1 ;
		RECT 47.525 150.785 47.765 151.135 ;
		LAYER M3 ;
		RECT 47.525 150.805 47.765 151.115 ;
		LAYER M2 ;
		RECT 47.525 154.385 47.765 155.255 ;
		LAYER M3 ;
		RECT 47.525 154.385 47.765 155.255 ;
		LAYER M1 ;
		RECT 47.525 166.560 47.765 166.600 ;
		LAYER M2 ;
		RECT 47.525 166.890 47.765 167.230 ;
		LAYER M1 ;
		RECT 47.525 166.870 47.765 167.250 ;
		LAYER M3 ;
		RECT 47.525 166.890 47.765 167.230 ;
		LAYER M1 ;
		RECT 47.525 167.520 47.765 167.560 ;
		LAYER M2 ;
		RECT 47.525 165.640 47.765 166.270 ;
		LAYER M3 ;
		RECT 47.525 165.640 47.765 166.270 ;
		LAYER M1 ;
		RECT 47.525 165.620 47.765 166.290 ;
		LAYER M2 ;
		RECT 47.525 163.840 47.765 165.330 ;
		LAYER M1 ;
		RECT 47.525 163.820 47.765 165.350 ;
		LAYER M2 ;
		RECT 47.525 170.470 47.765 172.800 ;
		LAYER M1 ;
		RECT 47.525 169.510 47.765 170.180 ;
		LAYER M1 ;
		RECT 47.525 169.200 47.765 169.240 ;
		LAYER M1 ;
		RECT 47.525 167.830 47.765 168.930 ;
		LAYER M2 ;
		RECT 47.525 167.850 47.765 168.910 ;
		LAYER M3 ;
		RECT 47.525 167.850 47.765 168.910 ;
		LAYER M1 ;
		RECT 47.525 170.450 47.765 172.820 ;
		LAYER M1 ;
		RECT 47.525 173.090 47.765 173.130 ;
		LAYER M2 ;
		RECT 47.525 169.530 47.765 170.160 ;
		LAYER M3 ;
		RECT 47.525 169.530 47.765 170.160 ;
		LAYER M3 ;
		RECT 47.525 170.470 47.765 172.800 ;
	END
	# End of OBS

END TS6N28HPMA256X64M4F

END LIBRARY
